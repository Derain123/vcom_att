`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="galaxsim"
`pragma protect encrypt_agent_info="https://www.x-epic.com"
`pragma protect key_keyowner="x-epic"
`pragma protect key_keyname="rsa-key1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
OLa2d+1qxOo4bCAfmAq8XLu3rNonHQ36hAEWR1hkw+cg2nd31GTW+PhvM3jDj8j2
KcDAFUzXTywe9hag29cDhrno6dDaiaQ1rtf/n//2y7iN9KxIodyUSjXR7OkqcCFV
QVJ09W6XZqNbJ0lH7RALbnmjeAI06s+OmN81S7hJfuG0VcI8FfDURXfgAeQbMrr7
vp4TSp+4RN4xHbyNecXu/RUKldW0cmTQnkJ2Fd8KmX8Wb/Q1FPQUDhmT+RXqkKbT
EoMWG65t9RVNghSUyr1cMzTUrsX2IICzdFGlS5ciJxyLgX1vzCQxeneo2YmyvxTX
Ty7uuoG47UWwLrkmu+f9XA==
`pragma protect key_keyowner="Xilinx"
`pragma protect key_keyname="xilinxt_2019_02"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
OkrznTFYwVGDdycUcIwq0iRq49Z4ogD3i+M7/vQSFLtGTeobB7VPzrOt1yZ8Pyes
TopKsPtGUfXTizXonyh7wl8NCyFm2oRQhJVuC5S4OHMTuTSwwrjsFY/8O+gtOjhI
UaEnnyhdiqaS4EbsQMFSkGmObnOm90MdxTi9cyDRHhu5XiWS8Xm8cO7b9cSdlIXB
n+03aYiNQHTD8q0xFwsoGw6mBIS24vXwjEZTnLHq3Vj4XPhDv5UA7UGJuGpyV1bX
/xJD1nvN/XPeHoWH3NyI8VbzUEozXsUrvpJjRbcuBUqakpo556J7NhZS/N/bnjlK
DAxpxOBTJSCaN11o7FRiBA==
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`pragma protect key_block
AcgLv28+/HBZV8k3cfjv2EXb/+dy5v2IwGt0pbqlHs7ki5wZxGDt0Fk1eNSuxLdO
/EhkFFTo+AV4cFYIxAuUQzMxkOsaduAtAHcShQxEPWCcTwIG5N+06ftgwdf5YfGn
vyzsdTH4H6zXIyjc4fEVW5j3W5jr+icx7BPjoHPRDKk=
`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
YfZB+G6bIkVOqln1purRzvD6J9+YZ/8fwpHP4LiMvyOwTP/uI2ebM22eyIb0TT1D
Orru/l4iQlTQfrGCfG7rUCCOuB4kaAGgCpEAYsIGAr8wpDVgxA4X5VRUpqV3+rpE
TxIIGhA/hONW3tPVp/AWG0QbbCzQv2Pi/4cwlRsLaWklpKnBHQ9k6e3YuDTJEyBM
UMXqr5cHPgAT/S9kVq9ZfVfpYEafsvf4wnQuKb5r4XMFHc3gaH6Yj5yPijIX/Uxl
GoTitIJf5RRFiUyNrx+VHYGfv3+W6vNxO5md2fNygPA6OpnBxY26b1u3jxY5V5BT
hC1DOhBlIsEhr8EWQohh3A==
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP15_1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
MoR135zVIy/8QyFCs9t9N3E4ADea9P9M/9g9D4M59/r8S31uyq/4bqx1XKmfkXFB
OJhnwN+Mn3Bm5KJo5vG263mgLQ0JZELdFqJ+cdgXKWmZL4TX/+hVP6Fkcag4gUhF
JOpbzu228fDZXkhus8EOS8lBoBy4GoBm7+rxMZJxK1679mLhYdfdXr6RPvuy7dnh
BST1VXQRw75jTmQEDz91gsCnJFdP8DBEBXzo7JTRLrCx6b4FXNt3Ph+ks3EBeKz+
81VvPJYMiAVdsRZVg9AlN4MpSxGNd/HykVEgnZ2WMIc5P3DyzdzunQGZyC0rTj/I
HuvLENS8txqNK0vjANe6ZQ==

`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 7968)
`pragma protect data_block
sCtZUQnM/pryqXNHe0V6cvdgbPBhbwUlSt4n7borovnUk2xZ4Ih6Fh+vSPEHLGAU
fGu/guZHpd6oUKLg5+QJLUllWxtqoYhEBHBMj4Qf/9ENJoRDGakXPErqOmb0r9a8
rNN3EepVgHykSCyl45zbiyIbszamd1edNz5/s0wNjhjawoqXPj0nynmRn/dq2yLj
ZqDn0piL4qLJvNDtTMwX7V/mu+X4yQCp/S3OzNHWDtQcVWmbJsGEfkuj43CT2exs
We95+dihlPrAfaTC2mMj0PIOHTXvWExJg6sRHW54kuaEtlFnuvB/fCMxZGhYTDmc
6Uk0k7lZERk4bb2vN3uCWuWbIKmef5XGDkNxGaI6Ysllqff1+p4+nQBqAMHDDhcI
dikvHrXOEZ/8DVnqorjoXkWOUw+nObZ7bXm/Ocn8rnxcg6bvr6oyU1fQmRWHEyeL
Fc9lJO9sazzB5bqGfP/81NwbKA3jOvWsyZGCGwXAx8+O9NB+bVn82cR9GNIiR3Th
DOkijcFQrltXnp0p4cjyjmx9ZnevqlPTBLXqiMkzDwB+Zev77sWmT1Q936+vYc1j
q6rgDyfMzUwvhgEaOTMdBIO2zW0eaM10JPL3rTy+KMe9s7zb19pCROR6VTymj0Cj
Et5l1xzPsgizijUs6KQrVOw4a7BphcycuR1VIz3suByn+/nvUoUcjRMZX5pEl9jv
TdgR79WPWvbrGxCgtBji4u2MfWNATVqBwvqr9Nm6LrcyFGgdHjPXJXbvcKM2kVuY
dyyr4UbXoBw4JdykpYMpP8sqgg61me7TrHclYzdACJll5hM9EHgcce+KLMoIkPml
DnhtVvsx4Tn/PIRGIjHGJWRFhCwxSW+Vx+IjLv0RCpI5siOJNaBO3ImJ7VP7hIXR
msAzdeb5RR/6z6vt1e1fL9/5+gtsZn2SSjtr8oVE6FKNs4gRECdbb4ZwJe8d4A5z
74ch925mMeaJPlO8ESUDeOSH5/cJDvrlJq0CH7Oqcgh2yaZkRE1eSF5MVYHlUEX/
zmIOoSQNfx2sXhY7FFYkBITIH4xPA2H+7d3aBZfrJF4EKeHeijXDpQm5I0YIIpO2
Nyuj5lCMJR6KVb7YDVlSgsGkK0u9akJcrg7YPBRGyDIFF7Xn7pajkvv+nfJDXlP+
ZzPiLch25u3YSssknejbxh9Z0Te0qqx9uu7h7FfTt5jcW8JqRMqrWSWs14Yhzvfv
YkOMgmbgqHoSPjUFqgF+DCKLPhLoWZpLRuIlYxKpI8vNzON5A1D3lY9g0XS2WhzJ
vbiNdVbLBQ3R5OdJwk32K79h0feHZWj5csyW3/s49ryerj/mwihLaQKubGW+CQ5b
3HvNuiPRBq5g4BxUHl6NU/DIfSQOVvG1yAXdBMpKj+WiPgL00C03GGapFZmkSeaV
H24Ana405LYue7NncRYinvMkmlvI6S5bByag5jADTT5shGYWiA6eZ9MXLPd6QTKL
wpb4UFD5oi2hHIFQj7FtVlbVdBh4GLwFKN2FzptfitQrXN5yW6PSre32IZ6gYwCO
wA9/kbF+/dTqyq6vJlckDc+PnBVVVfGQ24vbJ3iYBPSARFr5idBo5kYLtTeNHatB
8FzvPjkiPc2WfHR7tG5Vdcw9FANcOqr6CHfbGK0eYD82kYkUuMggHWgHM/pI4eZB
Kt2ZHXososZEF+Hzme79ZDQ9LJZPCY3Urj3UWIl83Zc+OxIPIVzclNfbtgN/sJ5V
zbXDZwsKsPMTy824NOp4kPowHH83y6JMcsmTRyEYUMV10YAj/ywaOLrEvu/dnFQv
N+erNRMEUqxjTX4LEYD0Qdxw3q9da1LsT8eDBDh6KwyyLjT+MCYiBxF+LCO+iERK
MQSsvH5cAYV9sywATus0WOD8SQiMAhS6QKMbM1jXS9F52iXQMMsAePN+ywKYgdin
m75aVjiVl/wxpGanBJ1o77peN6wOs5c515kmfX8VftULo88v41FdYlZs2KncFD4l
g355G9JhIPa4CiSprvxfoOVo6/FtoCGeGULvLvu5deqH01GkLcdBhw9YLqXQlMyB
5yyJBOwev0IRvnNtI9vPvt6RMuh1kv+pyB7v+lUMarIDh28xPbIweGfETlF/AL6u
WZjIEcTehFEEW2AmRqVL7AEXLLjf0XaXaXFK3aITkdit5+CUMK09BZR2Umvr+C4M
8piI6+2coAMGQpXpiXv3W+Nggze82P3VWS1ML8MUEMdS1HR/P7IbqefUkujtDEMa
1Ae4c7PQ/IgpOI94ps96HvkEc0Gm2FXcufkDDjLM5ol7ffA3bP6lE5CrMc58kEq7
6nTrQsUa+jv2gwvnw3yOcN6R+yII1FyVEe3J3I13BthaUOoi6yOupfdRdY04g+vP
qAkKv7UqxljBUHyUrjhU0SgZvtkrT3x43XDR48jPUxUGYqJJ9V/JBTCXRLneRC0y
rzgJC1cmegbKzSWdoFgkHefsMMSehM28aghWZ/DSBy+pj/Ux27fyGnuo4OdE+WXN
LyWTKsnhZpoxuu1RbBOzdFbtEOzeorIDpXSePC45jXcl2mLA0Frxdcv3YdqcWJAP
4XIuyp3ApJs8tTIqPL/7B69qg6mUKzwGMS9EsRsTCDYbd++b7yEf/MMO5kuEos5U
gzs7jdCQLFRWbbSeA6NOKy8GFm7b0lrr6qG9vlU/WWF7GIK6c1TdIkoMvjbBRlww
XiCDvKjZr36+T+eRsxBozap0Zka/AtF75w4IYcWkV2p3yMH34KrT/k/XIh+B9ChZ
//oLUDiTdHt3WbwYQOHZ8V3fkSGb0JWx80NxZSVPPU2+ghC0aHr524nqKJ/Ybvss
iWw9GI2Tx8sSB7rbrDLfvFrxbabQhjVHNwsR5sTvHFTkPxmzCm9IQfdWNyBam73u
72kkXbqsQR0fMuFVbizo783PWJkxnB4NotRxKkXn8bKMw3JZ/l2FEmye7Fifa3nm
KXKqEgM6d7C955A9IVnMHaqh8+rL0isSE8AvfaKEEZ5eqFmR8bAOIr+VHWzsxFY3
q/KGI91dmBKGdRdzHPNMwRatl2PdMEHElq/vrCjMZlpMlfShb8jsBbcQQzsWVd1W
OEBqEIUL6L/lr8yjV9f9PbnG4qkFVH0nfNVXwWQWXC1LYvTcShUPOXLj0Qb3EjYt
6By0s3L5nfZArKs1g9rjQbr9xoOa/cYle4bssvtvgZBi80d+DcdUuk/hXnn1i2z/
PoyJ/yspeYk0SOt1emXsAhUGwirlAIM8MjriBHYW9mA4p7p0WOyRWtVpFH8TrjuL
FCMeaFBtGe/Zdcxxe0xt517CkBM2KmJj+uk3EaIUmUeACHLWXcrRAfgZ+ylDas3J
ze6pDUFjDILzPc0KLUqF7HRN4bTP4iXneetyJDbWfdbwd7PzV/20W5x+F3xWiSTB
mhwczILfzScLvzG5Op3h+kJq31tj6l/XdvhkRMjGItQ3u+2SFOJNrfuqzzuLVBA6
sl7Hihjxe+8uSV+UGHhSd7yUgGDLWgrD/+eEijU4XD5gw71mXcnPrCBMso2ivvPe
yvGPnE2ZtUkW7+suushqc5cklgUGm7MZI4QK1SfAOBUQtRMSPr2WBfmhtYQ0QZam
T4XgcEpU516o/r2gizbIdoNm/sTcpz0p163lboEFmyRPR6ap7FibWS+lB9ycLmY1
5S4tTK4KVH62gEYxSmc3JNTISxDxZFmQJ4QITZCrEoyZ2Ir3T/EJPkXNsG00F5F2
XeCOhgTbAZAOHgSy1MZbt6EJ96BZxJ5XpAo83VDVLDHld5yLHoI/ClRVLRBk06FQ
QI2tDGChtU0/icRgYKBJZ2HJjMk5vHpBStOIVcsAQTk789PsRJ0UY9+2nCcvx9ZL
WlJcrsT6EvaOih5PRNBu4zV9HGNREi5KiDa8Mli5cCT9OUlFaw1+lpHFWdD/6qsy
rRk7V8pkhAi66c2hbE/s5IM/QKl0jh/7IbN3GMCRWBX2Pi9Hib1fmNC6lkWdUEQ2
YC1w/pmxLQ6AWjmFMNJqIaKpdX2P+Ly+I5FMg8ETiq+uCvMmpTiLqlItndobxxKR
EqLXWQ0TsnYcRcNl1ES6VB2dmIxDs1q33Qr1Zoajg1esy46KJ+9bxyTqsXnkCbto
5tBBxeDkgCV8eksT6dO7Q0rdo7+lfILr53sx/5Cs+6HgM6qNnXlf9boWdlfZEWWa
jOUbDAFfPIvawHpuE0aHfmmkSP+N6Z+P7vW/qU2ahpQ4/1ivsh1k/v8pwYlnJNnP
WK5jMa4z/3DFGWJLTI9WI2AzNaf6vH4Wut7Uot3vvKHS5cfwoHUOMz0H1d+5z1Sk
t1gU75jU2TNQ2JuqxvTiBCdS9A2rdxu7yA8Ut4H28RaDAqNWEXSlNzDI3/qxK4Ec
mNyMzgDlE1M2Si6LTH+R23kYmcaQ1/15cPdVFgYSyNJVMTXhVqgszLDNaKWHUsVg
B4lFuXG5/Rn6U/S5Dl6Hy274g/JYsR8nSg7NeCMqP4XSUZEnboQx+ZmBIy2akavt
iYwVWbYtzkHN+ceTCsfsFK2U2ydRteZfNE6dEtoFDcMCyRAv4hta8UUvzMRXU7Wl
iJ2UMPH7POwGJvNLYwP4UEWHGpzWVR+BtI+y5Q3pAWWgrkNNUijIE4EVy6Q3X0Mc
y8CBJQGQYFChuZ3Nn6ubmH5tlydLp430IIONhAnvQgTA6LQzlQ+htwl9WUrVuTqD
4fqdwRdyCbZoBbTlFIDecMpRlDILPUkeXuRpr3avsjBqOzpd7WC0bgDCwjumR4L3
H0bUnmygEwVKBkjMq0/i7j0DjJWSij9PTHXCbSF5EH5/Cw4sw6N4BwFoTXqO4xeR
eYF69/CGSFEifP+eOkl/Ga4xqK+89JBlXJZ25NRktjQlfe8hiBQWvQ0VcOPj2iMV
T2flHdXRj+CC6XXNGcmupWlj/VTrhzzXzeptaItlj1oWOX/ljXoqjr7jV3x4gWEA
30E+p7OCwPzlbIj922pD56wxHlgyZYZQ0VeVWfSrP3yo0dB4DeIWcaMaud1k9RTw
A9etle0HjFBRI2+QqNj7Eh2hFlb4FkQuleIHU4xh+Q0hDuWm4/9JVjTvuXftHEqM
bVfs6m+SddHypK338iSANhDmGgsYDx7PsYYsaarWe0m0jwmBSkKyutXYDleyQOm0
5H/VNAvOUi4giBYpOtLYZvdxBxXPJvKnBUFVR0pKdwt21BX/et+ITtQyWSJDCW2T
diAvHlZ9uYw3cgqIRaDB5x0WVa/N+CjX9ujkQ5NZYfmxRnhmqS/XBWHqc+1D+NXo
4Dm2imQw2RJ+vqklH4KeZ0Fe2YVEPqY2D1mky0M8ehitGhKpSNxnqyDMF+o3TsUx
JnGycgedpjXw4KVahM451YWfCstCNhOfKSQRbyU5vUuNoUqNzK+hKEkUmevw51zf
5pZCJg55RtA/R2a4ZKPv8RQMrpvBdW0d8WrHW5sLt7A+WX+4ZGLC8qYFktoDHkCy
ME/YtJl2OIbAppeP7iOeRU48LXGeKg39diJ++0/nfnLrsT+JLRkNLzTViaLfk40v
+xUU7P6uO7WZQUhsKNABOIunE1WPboND9a2/Mbs3Op1mZfSiq9N2LmazDvtQ7Mk0
2V0D4dSJ3e12iap9KZIqz7o/TlQ7BgrO1uZDS2JLKd/oWriooFlYxunYWiq+BajE
LdTEDJVtvaazedZNDEKlmqL7NpyLgLwAnGNQQm6ce3YQHgDhMwpqITZ2kz49+Fws
dJMgqLfDpoeEQcO8CYZOsbZvpKesy++inCKt6pqvBGHXhUF0cM4XIbOLJuGo4zrp
HUn752DW+bYJb+xYBkmVXAAppREsV6VeT3TUGV37lKsRNvfr9g7l89O9MetzJlRF
bS1RU/0F7pt+1RszADrrCo0QxG9HVLVmsPnbCjnhUxyk4of7hx8tNOMXtJwzDSZZ
95lhOM9vc0ZOiDGlwvsgEfYzzZE3LG5+MUwOzhryOKclWQDRZ60D0qzotsF+IGps
yhLPdtLHCS7bhC0nWS0ZrcvPRJ7DZrl5yQCDzU6yZNnBLIHWe26XXirXbJWtfOK3
2IWpqAhVpJXqXOFZ5zrlu+pG340nHZhV36SlnudLTM+te4pgWzOkm6xRn0SscCUJ
D+gX8WA+9Ycjf5jFQBDodBCyTKUxvhEP6ReQE9joQNYXl1GMJvWTQnz1A51VRtVp
3S74+Y446TW+TSiADzT1nHFgKOLwTXtKQp4IPgjKYb9s0fHt2oq0JAymJSoX257m
GCxTvORjkTdltJw+MJXt8SMJwNI8GIfLCaNWPuOd3TsXylA+BHadKOD0Og1ECpfL
81kODyGrfUpM2OOcD4ytat5kCULmNCZBvSNbgf0aacVowvob44rAuwpndtnIZymM
aRmK3iCinHxghDvxAkfuKRq1XZSiv2uRbLJwJDqeUoPP3z69hiJrpbckhKPbZ3Sb
cAj7iawQrKW/xt6F8BcjdT6nZD3OA8RaQoIQ2aDegDrknPrqQ0gcloGu2CBq1yfj
ByVzHp5aNV/DcrWDVJY9NayHcgTfGU1PZ4RWEp2ij24xJvXB8RiagK/Gsp+yALGQ
LRwYHeR3nAtAa32KJe1RbIRRjGgvIUrUVqfEz48FXeEfEWKKAo79duANkRu5oBox
GAkyCe4BrdFSUNAoroMGm3ZzRRRmYIEp6AZ7H7GfHqUzEgaOg5foNfEaotwd+QM2
yZ+7e7v98f+WTJW6I4hwrG1UhApYD+7Le+K3U40xfbL/ExARoiabg41rXOPYnukJ
va5skyLWJtXctn0Cwh1dufF8l5TauSXTPmJZSrnqrTkf47qdeEgZli/hST00JNO1
JcTF4zoatYP56aFy/lquFI3p7VuQqgm4UmxO0Ri7icaGYBoZOYAQ81ZjyNSWxSai
k01XEmG4WAZbyOCsawxDVCts1u9dy8RsjZAE0qN1zerGx1Or7Pb99ZpD+IxS8/kD
w70DL12uB6XbBYGVswP56314P727ygdMWrAI/c+HpVlpjxtdHZoY2YhBWzfFd/K5
TOMcVFQx6hQsKj9bklHWFJkC5JQvC4BKePzS7HDmxX3BJGCKI6nAid25pT1Vx6Vj
VQFcQMxTk5M7vzJ1oB2jW8/j4a6wq8jkvLfZKMHORVdW/1+u7fJ3NgPfPRC7GHOM
OtC5i3qWO4shvCBhegocvmtpnMcTxvfIGwsqTQ5HDKUTawVLGavq2rjdwjEm96uK
Bf4T/iD+SCAXTKpCdUkomtbBwuNaOEqQy3q/PJ62Dj9eCO8YMDU0TIXjV0GnxcOb
QI8B7zFi9alek/hjHEAOCnQkxbOYxOTpEtACpkF39Dm2S1IMeRZZVdKE6fAwdzz3
L1ccPv59JBZ7YmT/RMTpH6ikScdoPrChF40VvKyjVhT1K1XxvoJ4i2Arhis/Um5t
zBfUfYwclF7lnjp0m8GxoY17OFD65hmD3sqeZzqNvc6V7yZ46m8EIgjf/CZpGmyw
LQ9JitA0YB/F7uY3urnQ5Ez5RlDNtGE+fyUgGbHLCZjh2RwlG9vxI/KgrQcHgzFt
X9RoNP3VEUTen7GZin4+WaVXZKviQxN/1v+EmYZvQ+yteoLBi+PUaMc6J5FM6ws0
XV2exXPk8lVrPgxhsA0alA6658xUk1xiDKIYyTmruTO9vHykbwg2nlu3o/NHrwLE
2mQOsY6HVZHItRHUxhmjFAikys+WGGIRaozY2UBHi3dsli6PbOXrP2RD7N/QVXlv
XTX4Oagy4wUabFCYgG4wX0rhysPTLXotHH2hnymVVKQf+HayiAJq/o2lM5LrFz4O
FIXUvdKWDiQn4c+0AOnMcN/73+QV5BkK75rAwjPSmFvXDYPFg4GGVa4l7mVraTuq
UyyhmgJKCLkfesgB5qGppmhmBphsBbJSheAyC+0LYdQcCHnsgrvyR/79skvUKJWf
LrnEXqr+Krs9J2cHQH1WDwk7sJ3amrN5KS7Aoag32ZbSImPjhoh5l8yuwaHlxldM
NTRXuDg9qoT3mGHrih/qK2tDpYx5rIJga2mHOOpJZrqtFBL4eqDYxvsxV7+KGsM7
EBeljHZLq53jdVU46GAbu5bl8nUHHV1HmkZEm8pXV5C5T18SmrR80yJ9g3JHCL04
oQKx1cnjLxcXmAWO3zG5HRvkdQsLj7K1l47wkKo+E4HfJ9SHniqwT7vdu1PtCnEc
/6bqOgkE+yG/NFT/j9uH/DH9qemwWnZvRs//7gfOChRMM0zHgor0r6NCLkJSO3Ma
hTLTcfRVdQn5kgjIZqsmQVFnCT9J9jfrOjoLqKnuD/egKfMIqqbuWgah2gXXhwcM
kgrI4IPA9LBcpaO2xIXd3grX7kuI170W/LeMl/IQxZJ74+jnOxTaCKIGhShQ9O81
C7+dNhS7Plhg4w8fzKCiATHswAddeGN8Pbry0qx6JzKNF2JKvKfrkOjYYiQk5GG4
0/YFynmfRKSSr7/xgYwa2qKccYrDJNGtsCx4zhrG2kc/K7QgUGYA/GhM5BJVE8mL
RUZA5G7otgOhr2EWD/PUMJTfUBxtwq8p9a5M9zyAJ40iOFsUIGIJ7a6escFItf0o
HxHWYQb078wB7t9SzaS8m046CJQJf20Wttei6mWnz8V0X2+/JD3plyyFghWHVDW1
ZBhOOirqSU8IWRjH5yvFpcWZvMqEtc0Lzyb2dCIAW2ro+94yDjQbtxHHKe4o0NqC
+3t1pvJCCLaC1FfHiLEA6/ByyR8qMrbTg7of6iOiO8A24ibmZZRVJqYPclgEaU9E
Kwit/goZjVQgFcLRJYQBWW1MYrmOqVJ9okKp4LGW+vZC7T4YnbTJNxg20ELdcZQE
DQ81ldIT2DeK0FW5uRx8qACXlJWH5vn1tE80IB+Cu4Q/XuFZZ9/1NaSLY0SafZwI
JIah1EpnFbKF5nqiDph7ehDehT9XOyW4RDXZm1bETyRFdnOWP1ETQbUl8B8l1OwI
30jY4dULkI6yOAEIRp5VJsApmLOzZm9TeRKuNbYbOdvwqd2++MI6CJGb1JfyD91P
fd6E+7p2ExP/KVdp9rzfgisfdH5UH9jykzA5aFn+t6UZlZjmF5x7XqQDMd2kLRLK
w84msj0ZMMCW50CB7SNhoLfK6MgP5aq6QmAnkdCB+wdHWP5XST0RBKWJONX2YVXX
4fh4uVnextm9P7AgcyI4vU4uYVWU1ltVcm+4jFjLRXhQ8dWy3uNNKg2iiaGNu3mo
M8Yz1rjzEIl3xJEnaWwEYIxPQN/zAQk7tm0nil7kkqUibgDs5GBwcc9yzfFl2vgm
zZ8rBRb+0JsqoqOFDj2KI4cbWah+tLqQBKC31POjAHZkuonUJHqr47rwtZu++2gY
MOJPx6ZA5HaLnBRRn3XMwyarvlVK/wqPT/GQfq1R3RPoj76osJPZeq8RoC29nJTx
04O88895oBuIzqMyftuhZfHTZcFooPWcJdzg2p27N5kt+9YddFGBi8p6k8cHvNkY
CZAkg+naGFtrl2Y8L5ySAloTnMWW7Imm0ITi5+dFDTYvIZfWnpmv7lvPUiyJkjT/
PWaNd7++wmARWRNiFJMkzasnGCovXCB7psCzMSqcD6dCa5xRLZDsh/JQHFsamcxJ
dmKUeHFiolLTgUvijr/CqQB/IhVliaPPUN/5N9aq3df0eKn9Hfvv9ZUPm28gEgZR
IX7j0t2T5k9RXg/XzJP+H/LeUdd/OdxeMEzbYo1BDc17S5Nwk9CxTzHihwqLByCX
vDHJ3pJfuVKzsQBL11UAzknARsaWQPSmM2dH+Mi9vx6zkbD2VbDCfAq1wnMTvz4F
Sf0gHf7hdrxeDeP1Ij7RSvqSvEIB3dFIarXCQ3N6sT8dLhn6q7F9InH4e/IQU/S+
jQ68xRSOHHOOXhEPxLqwFAIukGQnhxFAkZXSe9533okpnkfOgN+ly9yhriSEnLYj
oD0MeuT0rbQRqWaFEImH/npShoawW18y/U3ABGfEzFOCrAypub0U7c1MItpIbLXH
eSIsRG3nAhS2c+6EYrH7HNVxBZ7ZRi4SXSL6RApLjnfds68CaF6axEznUJVEPskw
IO/1LBOneJB3vHriIIL5Rl6Qw6bhYD9BIf/iEIDGeINZVEQB++leHjh1b6QtdV+l
phcEPEfQFjIl+lg7+KWcl5a129eNcnRR/t6XYZyvFR31u+sysXUIpuem1NpPvEbm
RWUQuvIw/VA3czOszHPAW10cufCvQDgzPUrG+K28hEs5YUYRmZk/AwlADMwS31jQ
AtCNGfmPBK7ijfrFNOod0yo0EFnUFl0tKt3DZ+idNd5UU/fdTd+sRYHijoqZkP5D
orSe8WerYww9wUjSItcfD76XpvFivr6bX3lcySxBqJGISSXa3mdHbY7NdVkgJ8m/
p9fNyxTc8523h371bekQwjOfYPAFErs7ichEgJTC3T5n6H5M6VZQrUrtL+JqGQy9
KsSrOgrGKalbpNI2fkHOjgS1v1MtuNIKmp4X3Jjf5yeVlzh+y6ZcEFgJK8FbnAF3
CQNVIJ74imREzOuwmPS/wEwSUfDdZ0og5UtwWmL4TFvkZIm0zwR+HbwByVa8yh9E
djoNerkqKZT7oyL+ASFauOlyA3EK/sOdFgKtbj0rlvfzDZep51IaCGUaJl/L7O+V
kbrq8ew2F/IKrRibQeks6uroLrfAs9cSWNKBrgJxqSJ4Ot0e5VmDdVSNq/5rGYwi
`pragma protect end_protected
