`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="galaxsim"
`pragma protect encrypt_agent_info="https://www.x-epic.com"
`pragma protect key_keyowner="x-epic"
`pragma protect key_keyname="rsa-key1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
WnnxYTVvMVDuyEzy+hPDTUm2IPV147j865zYdcUaiaHvC7/vnUAInRcBJOuvV+1L
IBapwW1O6KkKl0wbEFlAlt4D0qclkng6di+l2BU4pyRaq4JMJPBxh5kKyR4AUgN3
CRSG0BrIG7C5aZmm6LngIS/9eO0Xaf4bDs8r/Tw+nhyBuEB7wD/CCUBK+hb6xiL5
BFlgX7iJIf7/BY/cmgKnDnvCf1Omjmava3+BD1YKXZiH+JI4/pH76vaiJtuMSCbj
rz7JTojQ1f2/ARasy7SHz6kqRrPlfcLKonNNMkCk72l1nCHx1DFZhQ9uJbR4gbH9
SNObrtbe0Tp9gV7bfctzzA==
`pragma protect key_keyowner="Xilinx"
`pragma protect key_keyname="xilinxt_2019_02"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
C4JIlNlczGESgECj5kBQIwQJl+ucS/iAzN+RLoqOutEBl1cqN+HX5vWc1R1uiWRe
xPLNQe4H63uGid86tf+Yy/TXXOrPwjYXaWK3FFKU3vm0vxmQy/TmQaHGb+33kDb+
fe7gUFxwXlSnHpOO2dxD+g0KWWfaZ5sMg5A2Tcrp/5xjQqPryFg2dyuy2hwZYvqV
i9GAN+kAHZH3ElBY/jHCL2IqRLuDvvbU+R2XAoyaNuYaf8uH6wmvJglsoqxx1X6g
z/EQiiznJA5vbnA279nDmbJcsbJN+ln6OzcwnxEnetlG8clGuQizMIVs5a1K5Hn2
d6nX5yfPHm31lCqGJ1qJkw==
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`pragma protect key_block
BUyfSxKeYhmR+nNy0wUG31ZnRGOeW6Thk8Dg5xoWcsbbHH7jQXYDYXpzoeUS/HOo
qNi5x/rdOrE5FSP7O9BLGzjNLkUd6m8rSCsPs6mSm3PEFsc3MSkB9S7oMe0yDUBv
WSYUK51bUwTlZeHAmFYPmMq7aSq4tO4ud48YSzafx/0=
`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
BFVMPOemq9kWujauMPh9cZzKF6s7uGIp+LOB/IeZ1fkKaUKMFT4QRRoK7Aw9TIeB
Hjch/pcoE4V5iKD/fS5LnhULxCDcUmRTkS7GIrADCLnYUM7BnPAXG3ABy/GvqxIG
X9trW7QbUAmfvuM7hNy4v/eQ4lVEKgdXd0JkWf1X9BhnsqHf0ge6lRVzpzC9JAIc
kKO2zB0Mh6AjpiFVnabXzi8c/xemhQSVLd3hbJW7ZTw0PqFkeGBL7+i0rD80SZFy
5ZD+ULFHeMCDTbOTmFJzLptD9OtOra1NjM7bucLb4o8pW+ERJjA2kORCXfWXeRV2
9NKdDCl4OsnmWLqpOC/cbA==
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP15_1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
u/W6hxwBztCDFu/L2iGxcxx4RcGRpjGLQuSiQlMwL4t717Sj9WTe5solVpOyxB9q
6AJm66OQEz4SBcKLEvkzcdq37J/CqJffeg8vlrMKVkykh1IgCxq0eGv3DT7pdByv
E2JkdXZw2CKXtGnKdHO2pV9mNpBqGJM7ypg1xny2/RUSxlvnasbpZilBVyBYcA03
A+ukHqkp79YjBQcDkIYQ7rCkBiUZwEYWY+vSm4UWtgjqiX7zJfclnvTRiVhwfBtq
A6yu/9v33i6vmPpK88wyUbF+MNTSSv9grrayOY7xNkZQ4o2kJw9lg2LDqi7kr1z7
2XijS8cQWXGrA6G1z25LLQ==

`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 8576)
`pragma protect data_block
N9QSZq7WjQNk+1YHzLRfZOkSoSyLng6RKDM+KQ8HbNLy6Qixar9CnVJgx1XmnQJo
2XzoBrExTCfGAbfz1vWUzufzixNulEzguVkGcc1JhUPjqPAv/JJQiyOLNDfbf7BX
Zynw/O7gSK1MC7EowrbajTIQvLW9BM+R1XbxjiIizWuVaCr7GYl6MxU4pFsC8zoD
VXRU9/ujcNAD56mYkS9P/sNGEZ1yDI1xVRl5ezIfNCPkbtmB4DI/7MJFi2M7WeS5
fprZjpvyuNEKIiOFp0khpuL/0R5Nk8g50OBfhE24TwvxTQxMP6pUJ489SbB8vLtX
BK5m3UNhgAzxe6HZft4ymo78Nnj8/Ry4rfiMzz/F+4L1q+d5BBDpHbgNQxq4jUz6
dnPBHjZTrXoa/5/asmEpR7qt6U08oxEzlqXqpdd4BgEmHPm2DcQ/Z+9x6XvnV6NG
Q1f/fSch3GbWatR3ohR7X1KVm/VjigGp9hsaOxy/vNC18qjp5K06ENFzL7wIb9to
e2i1iqN2CIGHhyDE8QA29mJhC4nZwmqrTG3+WY6Bfl2ora9WO7Cnf1B+Lt54C/ET
nQauTYLKBCkrMuAtTqSG1ZemO9Z+GELVcXJ4V4YMeUqNz8cNsMegxLrMmb3LWSRe
yuXwhvFi0fQjT+L54WigsRMW56exn3UNNluS+vjisRtHpbEuOvsh92akZxfynZgq
tre4zjTkdMpfJer+hyBreKTvyDI/71XMK8t1h9QNjKO4ebi8Uq0NMLpchmTauOh8
ZMzaJL/QF8pJQGy1YGGA8kIMIHrHSLk/NfB4rv1OtLywLsSwIw1N2LRcrWKxWadN
n9Vhluq6pfK09wHr9NtYPWYce0MmXdHlVNn5uwc2XfMpzI1mTHypn0SdQbWp4qUu
/ISCO+vsaIIryqpxr9967kEMEbe2D5926wR/vCrq02xGCAYX0W0CPCZRiLkvjUyz
XlLM6UHgx/CnybWtnIHBD/GXnLuzdtiZKpKS45tmH462KJjuyMsFY5S4hHHIHVtZ
ZeciBHzDzo0TDg/IoNV1b8jR7d7UcMIJLL7/j/mBjCxnUVwxKRj1Sim49bztH/BM
b5Mub5wG3CS2vyD+3SMKva2NSaPE/7yOXMWJuTvp0k92VX6CFmKfX42f+m4oryBh
SQ1RTW11TNORJurxXkWNdeyTJ1W9epchtJchMiMHx5H18yJU69rXUtDDtRwdW8WT
PLrSfVY4IOv+KVgtrQ3FO8qcbJbaj/9XoxsxPTo77/uHb1g8lmtQptSjZ6lEwnq9
/AGbZdmdz25MJe1FczwrkQiogMj6Ot7pGQ1bBNe35e0ERkYZjOV7gz8e29x4oTT9
5T7HF0sSkYjNq7vUePEhDBTX0v+Mecj6D+GvHujCUA9+CSuBxPJvCOL1+i1zzgw9
3SpHqAo7wGtwb/Rd55/hE2D0YeozrzQTjgSPRiwXu/TVDMs1m9Dhl6tFNUPXWs5W
uiK/aluFVrX68d2ARb0vooEgkvlIeSM+FiaaVcCNIxCzQPAiHDPfTO0Ds5z7ejOM
eKDfOOY3sNPkF3XvOt/7x7BBgmzqDAFgh7vhHCA3+KcznMm5x6SBqi1ZdUs1u9yU
3r7cZNSuVxosCrFxjIzxADSvaWzP0HKR7mFiGou98ndNgV7vIvCvyH8sFMNHeVGN
tCB7dpAuU2Qbp9O0qBt+nRpRniHEJODQX/iToCwgoRfwVE35ykQah059HNRfComl
a+WPvBjImvvQrVB0KazmCj+Dzuj434NQp0WWixCtavZvWqqM9htT+P1kmtOkV15H
clf/mQqPdsubS18kTMvuduUaxDEBAxW8a/cf9joeIGa0As0oMyKhW5tkpKl1LETY
VAOYuw5fZ5u67ZcF3XV6eQR+fJ07QHiJOJYTwJGe9O/CgnEUOKoR1HOZBeFHk51/
/U5cOjE3NjEjYdWDtNsF6kAHWpQm24ecchOtG7+st6F9ICtqbcX8DUBEW0EncDiM
X5lR4hUBz0ddHMYL6XkIh6b3vFcpwEX2PX4NNsW2s65fgqtyVgn+qqI5MjyQ7mUF
CSqcGZaQKQeq86qtCc16i79sUK0PrF84rCIIaHwO5mXjoszTAI8bVGxUxr+/kz+F
jfDu+1oyA/hssdlmWCylMNvV1yzzrCe+7zxZtCqLXlkEwdspltu4PkjCdGCveLK+
HM/sVznMif4rmqA2iwjo7Gv9brLUp8dExhCtaGoERPzTJ+n1RKM58cNxGfR240Vb
0zFYueN/10AgU+0qmYOGoacC9V2wefF5cg2ydiDQahVS8FZyjj0gvSxphu1J8p1d
HesGS1q1Z3Iond87xQng4IGYNLcG5rB0WG1q/uLKPRT1VXMC4EB1wbgfDMeNPtIh
e6mDavr2GP/Gly1GgZwizDRtNax6JnS2POLhfAnF7/Ftoe4gNyiwLASzZiCV5ts2
MPDrH0EK0S05yOajEUp/+7ypRcae7lkqZV0vpy+1CjgFZ0YkwkZqu7uwTBwXhggn
+ri1kWveoCw42l1Z/dWE8R6r2C9EtqhDhKf0ewsvzUXiLuCPOzty6EgNBEnPgNqv
OmTwpFPh/dWLRwGXTpWKcus2HyKHtC+x/epMftMRWbZX1WjU8Y9lA4OF3829xM1P
tD9fH8IFVyeUCp0mV0tx0uNLEqJ5OHMGyKfNU49pMdryinL+UxMOPL9K1RMJI3Jp
SdJJ2eycVkYtNdzISaIRYEajo5CxEIWfz7zujJv1tYvlqTUu8eDg3CUpvI7R1yRX
G3pSbvEuWh7F1o+TuyiUNmdKpPhGsCvagL8vmyqbe+mIh7ol1i5kS2JnRt4idRaq
NI5bOB0ZZPJpeuB3vzsBUPGTkaBuePv38TAIKfJtY+s453Pa97sS2GATpKpdAK4+
9MgzKGpv+WdB1DMOffdvmFJcvyb0EB8je7nk1Ec6RXkx3hYmCB6b3vTVRqiIqNvH
UWm6yb9XCST48/eM63c2mUF5NbgA4rLS3TDKqa25ALTpGHY9b2vx2mDmBWGAWHCY
KpqrAUBb2tbYNNjacLeZ/RvY9cuKpeptoqZ5ehWRRMw3As+CKLqnQPdsqw6dkVl2
J3QuHYusqcqFOFeBpay4ui2rbw1X0ikrdpj8970oksaaNGRpbXitlHPkoc6uzz07
KyM2rTZYcc4Heg9p0Klem0z7UjzeQ4ndGUde1cG2JQK4Q+aQ7h/0CvORVSSW717j
sAoFFoyzCi0i/atqjiqg+EKQC5i+0rYji7fTBkLgqFvbtxP9t7B2is9sVGUFmWiC
LFcDsAiRFeDdE1BJ/eVP3QHMNoNrleqz2tZ1giJ8CEXI31wzn7suknsDT2OS/ctU
cLvJaA92r7gN67wgJshFse1lp1XjBXhMI+MPiXHG/Mwihm/Z9r5HxsGLrkHUD6y8
uKgqKmPgtiErXhEO7NLOOOc9+bKT72cCYoxpelY3vywi6OccD3QKEUN8Co7i8soe
/Xlb2Rnz7rreDDj+oG7GDxbbg4/Uo30VU/vPMHwOU7Vo5Mzp/FGU3eHZx86FuynT
6SPZu7ePRVzztHsH9xqxkMUK9NGTeYsGeWnZbxDpL3psa9HcyRpvtH4ev27FXSYy
N0bp6MUMZq2OGEHp+5LYNTqPbHzzq0GPshzW7gzTVPBXCKcbpZSB+QZXO5IrO0Kh
2CFYsVDc1XBT9B2LTuOPD751B/ZLl/IgBzlEG8MrlNXEKwDGf+nl9i0bMPVKrKKY
kb9PPkO46qSMdk4faTsKpQ490/60n1oluyABQKhu6EYKk73J0Fs0QBrupyczcOaf
yYkee9BwNcvI8U8Xizh3mSILnZNlf0I7Ail1F8do8FeAcjD4Cl/1F2OZuAXzNT+v
YnoKvWGGAswIo7brQ5gBDRf1OPcx33gC3P7ZQFx7zsVtfPFv4GZFUY+4X89/ncTf
TAt7iHpjYeGKBuOewAzh0hEsmL5B1n8pscMsr4dmVuS3oOwy295ai4TL8WEM4XSZ
f7CvFoiWKYwjPg6w/JzBKdihdxQk/SY1H7K0J6a2YJJ5DojJhQvfwSU41sCmnBor
d1FtECvOBrktN0LSF4xKERR7wPhsJWWQKdCKOfLFsJE+gRjyvcXeYe61MzTv5OiV
kXPX134qgeRaCeXEZSrIz2HidiyKocLvvSL54vQUw0MCHZutC75MoW86H/dX0LyK
nqxrkRpJM0CWydWiAlJRaVaKwgNP/1p7zd6Bsu2bBhao3Xs90cwzN1tnJYD6ZZQG
qwNWNXQAfXvpZQ26TK1aN74dlnSah+O3aOMA13PFv4hrpoJOUpykBPW/5E/dgwjm
KD5qLoIf8vZaLw5jodnNqqYOIUPqrBTVf3Pgb5ee2dPGhTvYkKtqp2PUo7Izv9Vg
ollAj0qdVSk1axz8fCgXBCNI4ES2At+1PdRzMgIKudexZtafJJBKC9WzloRzYPnV
eU1wD2JH21IQoyUpuf0FrJ8KYhXYIaUkEWtbw5U/+KjlQZuTxrVlfguHW6+1djyZ
NvnzAC071tozsAO39QFoWHmTAtQitGVwrFEpAK3VPFlxm6kFZxnIz+djjTRl9T3g
9NT9hRwp2ocp6qDSxYH3GtR6XfgYAHV6VRYXMq5zlG4qwM7mfRUXWh1Uny5YLidQ
ux+1y8FpnFDrlnE4IzCHi3QnaklPuAXPxi33IioSSNGtPXOh87tL0wRRje7tm7u+
ypeXhE4tnIqYDFHLwhbETp7rchZ/LNvqL5qGplnbwQtFGN2TFXyIlHU0tywlpU6Z
NNMHQ3dOOFIx09tHoq8hsYnxAVSUYBEFgauyEskhJBlem0er9DnSL+UwYB0CMUeX
HcycmUtd4sDZbI4pmxg9LWmtjDjyxXSYrMxIeP+bc8DjinchdpfVS+wy0tZ425KB
g7We4EibFh810L8LI5ADR9CkgdSTCJG3EuIdf3XUhcIB2olV1eB2cXG8LixgtdR1
PnQeMHIFi0MNhD4V0uoSs5frlTU+BflKgf2aTop0vtLkjI90reXi4kNnij+bBL/P
+RdXPLYYay4vYE/8SwQD1kojubG+H7+18MuzpJVr+3zEhuqsf39R3z1iujJFJfus
XfXshw6nngifMX/QiU3NiqqILcBtp6PIaYfBBFAF2gla7oi06/gjabvl4r09m5zT
7fMXvZ88YqyZIbE2UMLfocoV63+ykUkpXtMdaj6YDaC8EI6o7XWhSNohh3WjuwL1
+DABKQ67INBZHTi5T2ezMieJb26TwOIUlVtm+1zkBZHolD9twEbgu5DgVeDfgJEJ
/N+lqnT1HVckoVoq5aZVOcy9CT4GABVu+nvt/jbowRBiMVCS5Bb4WRn7WtpLwNzS
B83ikyRV60bWkvCHg9teQDpdtsvroheKIh/ujLmdZdO+4fB1G8JAJaUN4JVsA5nf
EzKZonCnuUj0pAFL50xSh1Nr/uJorI+BLQSiGlabudvotLukykkvTMuYc3trJOAl
O7LofvH/jFEAEj7iQC61ajM5vImQGm3ZoP4iyrUN3CdG53MEo7Dt+MNRf5sd9GSB
2kS+NHr0VGLSpv2Ne27H/YwpD3BmRIz+BuX+55sGIFKV62gTGxbxLF+4pYvX9ysr
C0ZB9e+RCTyb0V180nysFcTa6JESnhPsjymAum5y/PtQNus+90VBeBg8b+Ao9L3c
JJNaUTDdXCE3xwr66dJociEKhxyjjLL/0SaKCIexavNQRu12bxnG+U5pfBezkPLr
ABA0FACq+/8R5xotuflXVibuYvqIWGd2+3L4Hp+MVlFAjnaXzKOsLxligwix6DLJ
6ZD5qnkE+ETWKURQHkKAmbtS5xMLF1PfasD6sh9ABsGV6ZuuCrCk0xcdDDRdLsLr
gCP9Z01P6GLFqigpuvWVMxleQlii2YLFiOEllGPYvlM4zIwcVwhIqWEnI04GMGZq
1U4EFL6V5FLPZ12qR7QnKjPD96bCsiwLsVzK9zbvDvq2LEOn+dm9FZPPGKW8WGWT
9r5TvbOH9ZlvU9ieZ/Oy+XIPefiTUHJLDp0TsXAUq282VUSK3EP6QacyMOD1qjOs
Nrrz391tqzOfGvPhtWQ+8Gs6Nh6qJNMl1qclVfxT225atv36KrZobzVGJkP1Se9W
PCP1ozXc82e6YhBItLaamS8grPm5Sab+d36Uw/UzdF3GNgKhi5eOlOeVfO7XnyfC
HARdjs9tNYKr2X1rt+XIA6zgib0RayDgB0D8ejNSHkqVVyu5DJsJttf2hIEpzE3t
A0TvXnMk4pRqCkGSEhrwt6Neh1mnk7VmZJbD8nZUywO+kyRZrsyZCLSfwVBDmykH
9P8UnJviWauDeORsQC2ALvJ+axxbVvhkepoBnFQboI+XCjFK0GZ2RggXZ2ZldAY2
YbgdS2pRlHyiOlSdvYwhIvJIPyLCrElAY98TBlBZz0rb7Qc1CAWqVWgTJXiWWW45
cfLOTqBZ4WIQRMtkyCT21JIwtNmCTe9klpd9nsH2G/nebyzLvlZit1hKzA1Styd2
iv8dEDsmM1ZcMqszVwdzCPXnUhptexLW/YVDYlxW5vTHGVJlrg/zOE8k/uMwH8A9
RYHNClcsSpfNQ7ixhN9eMAPjIn6ZS0hVeE1L2r9yBTVk1xpbY/s7s4lL6XkHzxSY
kf7f51dNEQZlCxkTuVMLp4urNGcHvrDFQ3Ds5NqKfXOnMS4BVReDWrql5qR6Ue/w
kWQt94rDvQAY/qad63tB8KQBFkQ+A1rGmu34jGF+SLM6wsk8TPZt/aofK7iVFmi7
h7bv1UOO8lsvQ2J66pcG/cYsouZIMicxz+vfF/nJMqZ+ERvHhxcTv9UuwDrqn6Dj
3rDqcV3PlGB0sw5+dG4DJwu7QQ/iAqyKUHT3uZS752rewFZYPrp5j99hxa/TfB9s
sytq/oKSJURf2N1UEVQ0Fiki9ULi9IQtG4xqwMSF8RvPT/1mgPFz0lfRjotE38tK
QzToFkOjbsJ1oggoDVHmvdRB/bCkuMbIOMziJv543nm4ckfRcDe80Ic690+l7DGV
yJZfSKAvopulS12LqfEf63ORrneL5OwPRJBrWU0CTfYZ0MmbBcxtt45OPyFPDA8I
nbre2y6dE0n/R4NjGjDOo+jZI9jpr3B1mBdF58F5eFZJMCjx8OVHBTNY92EBKYuJ
PoY7xLH74/c/qx7KCGVpnYjVe50lb/SWnhYjQC6vvMGTMRCpbjOWtQzgUM4TDZC3
yqqv7nVPvYLIjvmNdMQDqRvg9ov6c0iVZw4SfgUbktZmJuhvolarS79MtaxZAe+J
4+kawXucqIDhRL3RdEHScqMr+ch+bZ+6KXYKLyupzxZEc7rzXRJkAu8iLUCJaOgv
g2N9w1z3f768BXxFWPMvcj1QzdZ9x5ICW2+/eS0kZyaETmM7uiA1DcdNlb/h/tyF
XcWzTgJZdhyadHSKcMggBY5rDV98tWEaI/8AsnyjBapQ19O+PZosdGuSuXwCIvzK
YkrM4d79qgKzuDyZZpMbxlzM0lFr2eQ5UipDlDVReHWGLjhaXYIeIJLnMRA6t3zY
IPRnxwD1VIj4HzqU+64lCFSS677UVxG3MLhpGrOatYA1bwfizah72lbVNhQ2LM7i
nEtxjffdplHqzonaHeYPFUDJ6VpAkrBr54z/qzysSfeczQjbJE6TU2J1AZF3hpUN
HDNxEm3LwCcP7pMFk8fZSrfc4qlQNvYib9tQPN+Tq/GVV7FD8NCw9jRCTB1gXlXy
tw1MLmFAg7c/bgcq3bR/6z4a3Qx1jxTZPDWTvamJQxd7MW572WNlSGeHvAY3hdTD
Ajc7AX1wuh3kKjdGvOEadg3Kar6c+0pdn2ryPNHYg1cIV5LL5PDcluTJ7lABCsWL
aEvayGCmlBWztTEScEThHTg508HXJLPvXTYAL42ws9X6Hu6ak+d9tbzYM6LhQL7Y
15opMyk9dZfaz/1sIr9f/Iit89gsjoKb4IXoqwh2EY3GV46MB+FsVJg+e4oXLOQS
XlzSNwdUmo0+WwTCm7r0aYiK5nLUJ+vXCa6Ezlt+8pwaovsMNK7u59Hj0t/0Gdf/
ZPjoiKuvvdYm3MTZuf2WC8QQzifzcSH7S2z567eZuC581vmCLBKAgI1YfURL4fta
DKc5l5B+dsrbZibr7PdFDw8NfR93FV39LEsqsI05bfENhYLykwXRloOaTpw72J0e
dlBiEWqFNHWw1ABXYPqFONy5L6aCRHpE548xqjfyiwcDRM8pAwPQ3LAcymk6poEV
V5k1qlhDyFhBS4oVnBzX2CF8m2AzA6yZdBA2JCxDuIEwwVh8XbrLDL2x2CjBhXco
o150Rq32qBkjWdCHod9aSKNxp5DtzMNYMDjjJp7wmsdANfIAywsb4ubzguMmPWtJ
+5I5QEpGovcWGyk50hsW3ApKFztYM5HUFNK0muaaPh1fZm14x3obMQWh5xFP+KiS
z7yhIEXsCOsRtl2BG57Gteymx0dm+Ys/4hF8J8L93CuxdRZL1iE16dbM5yCSDO9L
KDdWUnhJOxs6mjQBODA19a5SVNMT5nSzJhsURs25actVl5pwFBY5KSyaorfVgt4l
owTzyrYZWprGTD1eo8F27LQsoiy/M+t5oSllweHwm9VO1raTnH9Sbo53MP8XJ/3Z
1oxS0+2V2ErBjtzZAtMMREbXD/2MwBw8zSJseGqjnCUaMym2JC/9hothHJXJ9/7Y
ImLWXx6vJmJejbsGiwJ41w4slcyyfejSrwAwtv553xyijZwkYHPSq7v8zT03wluy
nKPLtLpRKTssJj7FY44ncygFWDxSZqonVKFZ2Fb+AT8szlPDi7IG+OBHOVoAXknS
jH/OVDXGaWiJX1lJiroigBANbR2V11Q5y+l+8B5DjxyWshEoc23WnYtTStgl3Nl7
wsYhM5jAXomS+XwuoRVvi6l7LpM1gRyBTzhxUmeKSSDgSeErz8mQa31RBAqmmQmE
gV90yi1kb22B9va4MRfKGX3ODJk//KaLVteKg9hg84zksBuFGyzHqsqVNKvbbvmC
9WT61E7+KB0QMnOBckM+Z5exlVrBl7aJLaXhIXWfzuZ5xUW2tmcDHiUb/EsA4Hl9
HRT4MA2Xgm5jQtLOt8CMIVKNfjZBCka1pNwo/mpT+j2pw8Vv20bkfkmlvepQAMsw
aCGqQIFYosfZrzzxxmedUJ+0/d0yyosr85+Xm1fL5bXxH3AAN7It28Q6em/VzKlE
ZQHmLUDA0eAy2KscT/YRv79NW0J8xXfetZSC1bTvkSCtJf6dHOOVTbjqTiqidpVo
tKylTMEZJJQ50qyB1BClLfgZ+l/dB/JAmgBW/qjepzVjLyH2IWOdSvr3/Bos5N5Y
ykomkHrtsG3OQDqgQd+zxzPLI4o5ruxqwV6KxA5Cj/TYGpAO9BaEMHfgfFr8hiKl
4RIgvRNzC20traijXozp/WOeV0dlvmJNTz7PLYqUnxaGHqd2PIGpXJ4MlMClLgwc
J1q+YFrkysLB8DU3uYL9BKMkDp4Qqj7dcfB2DWhMaYznnneI3MN853aJ9WHho8rW
Ftp7Ow5jGxt/kCU/TxTZ/YaEyJToiQHtX/DaRRv9dej11fO+RR25gO1X1xyDwzMR
jPRY/HwdaTdPPAMYLVzQ7rrgMhpGyCnkW+rU8sg2/8xd6xcZTbzlrXzpndnNXDZE
GLO16EfLLMtYe13uCCGSHGAeQeiI4ApphdJo+mmRitn0zVWYBuwpKjMY1qNBgF6S
9d6F/Tq4NzTlvstYUjB9SusvShuBXfnU7GNtL7rGenuQcFFepjc3x7uOV4o5TgpG
Ynk4pwvyVYiD3azDPd8/ghbG8hD5Okaka/s/tMB0eULCS31ZdtPnhq9wsjWjQ0Cg
RXVakTS4tqFKsNNESiBHXzajzO7NKeUuAhLLKlQkUhydC7x3SUuALWYkpreZFdFv
hxrFtb+aN/DW7qftszZPf6Hk1EAcKaHhqguUHG2K8ic2jQuOoOLEmZt3zuifFLrr
ESDRcKy2mvlqLWJqDo2TqmB31OPE8nJGTAnjCPI/NvGuDWctubVD7FfgpYBnZRH9
/k4Qjqfg+Nn0wOUHmxXbn0y9L85Ruzxq0bx3JamAALBQVWWYJwMQzRkQC8OhVxnz
54mxf58Dw7I375UFydcTOOeUpXByqKgmUQuJUUo0rXA99Xu6zGE/bHQ5vvYJs0xs
2KEOsSQamJI3ku4Xj8DcZGqOIBFo+f0qzLEHn5EXXQLY+w+RxtzBlcGoVTVHYYCW
Q8E80XsGoRt26fV9eUC4Ea5oycT9NBPLY9zYyo/uKIonHdDhvzq0e0WmTycXW3WK
hlNktVpBa/Sg4MikS68on9NC3Ztgp2PWsKLDwwR135lTnSPmHFRR6HoCojZ4zPFF
8THreEWqW9eQmsxC4YWuyTxPxOJbnT+vVk5ESvJOWalu+f5/HZGD7lvSN2obYFow
GYePkvr/UGeYQB0OE+LC/4lPw0SlFWRMDbZACkWwQqk4h1/y6NKmCo9VtWPSHe+5
EOyh+LBrZHEohqDdC1VelNug+v5AuW3dwruqOWjpNP3owlU0GyT/b8B/Yh11tCit
Zwhu+osPZ9XTJ5zD83CuYwdOIR7Ucp+JdDsUeFWqQt7gwq9vnqRSqUmdvHOsRup5
AIhXQnSJqKgPvccKoOKJy9+bXMeOiV5DIeZOBc+qycX4snP4eghJwpvvaZCl6Gkp
65LHHNi3QmLace2B/qPqobv8NJRIDgQziu5v+JIgJBr6sZlEO3R1qzKFKFvKK+V2
rWf1b5DBhpj11tRXLYCfIeFbGkB8lCeqY9fVZxIl2OAa+35iXzMo7Xvtgrt9sW33
c8XEqsyoIvqZUggeuRFdHVSoMFnaAz910Q2xkT17gY+2nj+oEVr7xY8XwcB3/4E0
UrI0LIN4NcEgz1NEvtwbRF6hTWkmaacGYOPHpC4LASw6U1R27zax+qWHQC4RSsPq
Ey6QeCq6QsnQf5Ei1zS0q41EzKTNY12nAi7MFrwU9DjbsgVajXXyVceDT1MuyRBX
dvU1gI5kJU9SRvp45NyHazUMjsUjhISB+FNHBB4c9FONaelFTMeLDaPDDGb2USvJ
za3+W8cfCD+JRHV5AIRO1tcGv2C4HxdvGAFnBS9Eq7jDZHXogkpfza2qshxvUwFc
N1sXN6O96sF71+gDpYDbMsFfQkiMvtjLH+kOLwOX3iLCUmXiWjPvGwcq3VvlLx+e
t++XlUoM8LMqqTPaP1TkP7H0/2O5m3kJq960c2P4+rpXOwO9D+w4x1trROFctfEH
M3YQ3U5etqyGvYzCHhezqCM/HwZ2SofQNIbfPE8OoV6pz0cnM0ERX/H5di1t5NYH
TD/0pgUHnaCcB1ktnRgCSPOIOyZrQG/a9jsVLlgVyWqT9F5vztoe7HZ/jCrfHblJ
WBiV6W1+amaCNp1h9qUQUIQzLPGbpRLOKFge7hwhqYKUBOezTpmC6PShoC58hnwx
SjC18+0wJQwZdpWd2S8ruHvBSKNb7n8aNtCkSDr4aCk=
`pragma protect end_protected
