`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="galaxsim"
`pragma protect encrypt_agent_info="https://www.x-epic.com"
`pragma protect key_keyowner="x-epic"
`pragma protect key_keyname="rsa-key1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
WIE03sbUNr6z0SS7xk/gx38FS3PmisFnBoEEJDQ6Iaypgmg8KZ5A7MUZGz7qUkCl
2h6WwTehnaqJAWuX4zuy4v+ydn0EinZGw91xfJ3I61mUDVInc9zVw3oLOvzeB66a
gWIQQ3e/mIuP/crQpHm2lKonWQL1wtvUQ9bGhBd2lQ69yZECzgB5PffQouLeRWzX
GIy7b2Zu7x/ffjdxBqja4txSnMglgSuVpiClWgYd3IvTUYClMHOceMPIjL1642sA
oE+VbqJtRvO+MRKXxHZjO3D1l7AfmUoSkoQPb+MkJxRiPnXn0b2SQT2xTnfu9N2m
Qn4T9xrTsmU2dVq7MyN+OQ==
`pragma protect key_keyowner="Xilinx"
`pragma protect key_keyname="xilinxt_2019_02"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
oPOdepAaSow4IqvfNS/LVNM3gdRXMV1282nBTD18fcioyN2YRE0jCLwUp9xV3uuz
y9wtmwyK+CE0PUxRtyAFjpcs6t+3dhOSUzrbkCbb38qjfMsTa87ATVDF8b9ZeAnB
UACRb5vOjRSLpEmWcl9QEmUxVWpgeqyP52Xs1p3FNwFqg9uix0lxTuC7+jnbXUJZ
EYUM6tZwlI9bxTINY48LTKpEN0KyZuTsr7FUqSVnRJx/e1CG8dxR/MzNZpi/et15
Lu5RQIktweffe+HItoKbvigWdQWKuc6GK4Xe7Z4ARd0E6MkpYUOwTH5I8TJmHJgp
11Asd7XB+xi5iOCJC8JP6w==
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`pragma protect key_block
IERI91aZBl3QS7mpiYUTgVcgrjm2SiouIvK8JXmdLo73BksKlmlGT7A9mP5RL0Rx
2NNYHmNP96F8ZArkmXDotjaJyRSdfLdW0mvNG68eW0cgjOXlGpc8sYE5oQEnhvnv
GW4E07z8m+72dlA6JzRPCOHq7eUvgmnOPdcfHcDHfug=
`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
Wxw6j6zjtynN9PWCexce+O/cF62nJykqvf3IUWne7Bq8lXFX01doQJClHU/KyLqr
MOo+0K01gsPwEEquBAGzCpnDAK1tIsOdw/nm7uubEL/5YBsXOcWTS505k+bM6Ev3
CMryK1iSNafYoI52bPtTSq8emxarwY4fiAfF79Ed3EQ8/rUS1BL+lOruplI4iY2R
kCXAuXpB3yEEN9/UjAqsIAzlZImWviiqUsg02nSwqhlUO4OGBuuTF+1oKgvCNHLW
wpLuCPAIvbSzpkb3x5cn9sPVhsEnLNp4rVRB/liEnxOpFo1uz6Ivbe0Yk2JGyq1a
63SU6XxBnUaDYQ3EJ3Ya7g==
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP15_1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
UrcaoZh4gBLt32/LjhHH8NsbPnYLuXYuQqCsBV3851Lo+uoAczzKhMsd0F1eDlmk
7ftfhCxOE+yNU6CjaJFxH+IgS1WRj/mlpFamyA5DJkGeRynVU/RNALmYWLfkpS/y
gnGMB3oxcc08zTFVnxQ7cWRfx5dUbZsBMwxog7gtU5sG1Q0sPHuTjH/ycDY4xW21
KPKTMLMDUIC2DLJK3Msys7Q8PWY76A+uRmOL6Kf0Ii4KJ8gFvJjTHq9nNmjbROPu
iB5yPvsACt/qO8mXPfTmRVVMYUAIfzQI7R4ODkML4/RfoSTnGvej/aeY4SOqERWD
e0yDRWJ8MxPbKIWQ7J8O5w==

`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 8176)
`pragma protect data_block
IUyHKlniirs1CM9FBIk7JRtN26IDMOD8vCiR4BlYAD6B2MrfxEBIGyOwqQxtdqxe
lCBiP+2/di+1m7mGlGzLIe8piDmhlj1AsksZRCwMTkZtZya1DXpUbgrVqCZIxVW2
SvkUNEtwNcbXkDtNupr3pnn/BbSWKlduE8tlfwl6DJ5by3H/O+/xUv3b865/RQnB
fe6yTLJYCp3uHhNPUBfl78kbYR08mHlBs11VjmkK/OAiMqhusDP0++hCsbHqW2oW
sdEC2dSMw5Fy3pNorQB2zS7U1Nkly2orskTkXhKcR97jfmeIgZ0oijyq6whCRSgt
98MezpgbMaZyRelnE1Kil9t4coVySM1m8RAVXnZXbhjWUT4uEe5At159lrYVP0ef
NEAc9+uZEiN+5L4N/YoNBlI2aourjY1noFZlUI0VP0pqCl9PgKjSOtP+fn6PtClK
Up2e/tG6W1Sbz+nl3Z3B8CSCSaBDTsULnOxMx7Goy24Up1gdIdG6Z+xKdSB6dGE2
+m08j4CCu0KQV+U3Ld3J0QQXnojk1g4mZhc4dv9nWhcNBOyB8e8D5c/eO6r266rU
YY5WYw7pT/qLpme4p8Gqrptx8+kN8cDkG9DWJb72D4vh4hAXFXYbU87dEKI6AM4x
Ij1sSTHXiCijpD8ndr4yeSWlZ7aahwoMgRmy9U45XcT8c339/8cAtdEmxJMXYh75
A6+k1Xz5OyyvUAINUGccTYseKF/a2Im3vnux2Z80IH5RVSaf6uIr7q0arGJcpamq
Fb/9qJV7VprMDcGdeMXBn/NI8CWEV19bggqIp9t8LeC698UDMMj+QueyQHd1VZ7g
iaUrDIsSNZM0oYbZhQ51SPVFfRIzOzM+H/D+nzs3eB8LJkkvsRnNi6wttaSrtK9K
muftxrt43yd1cMHqK3SlnACfqBUS9/EhL+gzPannR1O2cNhHPBRtu7qxV1CxIp6g
ZmdR3vLTCTUrWLhovD9t2jpXa7Fb+VquLFIm/yRr4FdD0pkua9YedjgiPbI1GAEJ
k6dOUMEflcJ/waL0mvs4i0avoX0TDy12rM7wmLJTP0UErbmQb72LJ8wT0ZLaMKAK
ocIdtP3dwIWpphiguDxuN2dP+DwVQ6v2TcCP3B0/YOxkoSxfjHJDzSx63yofTcXM
OyT097q7/qBXoeHJaEhmreKEsWakOV9UntxRvJ8gvmCP433y1+uNXG6OJsQ9ETlj
wWRbt/2NoG6n9QvVCtRA0xP7OOjTLd6mzYjdWVU5mc1CVTTOUEsZkp4OV+ZK+Ms6
cyI59iPxfdjUCvmvbcr0HORvM0CZofTpWsmbmwrYuG8n5NA2FSQcTgwJ9KQoOWw1
HppFqf7TItZHdn2gWv2j7ToPSnpzHBesvlj9/bBOXxmVVpOgeP/AKjBhpY9P9z27
avEqd37Pq62hf/fp3/it/kPClf26x7qMsKcHnt/0xWh8LjZ+NhLVqvbMk+nQjnST
cgu7RcXoXmDvXpSeVY+1qmH48HzKwFTvtwdBwLcsHI2FjW6Js2sVzcyxqnuD1Wzw
TKARphAiK1V26Bi3pXq8sGZxziU5vk8q/CUs5mCCPDJRVR3OdXn2HU3/bXuWv43F
D3HR0J/op8uxQcmKwvIE2ekT2HZLUThm5uuwJvTOynRkd56Knqwlb0umIQOoJ2HD
h5kINBytLv8XgXshupi8L5MyHkgPbscvCu5+CaOXFuNBkXiRtRLJ1JwL8OjuCaIA
Nb94Isgi2tKqU9RB66Y4W4Xk3p5M9DjQVd4G3OC72w3ZQC6gY3V6uecwvhZDrbJZ
KRxUoPEPD6wABkEMZj+BK58tQuc3FoddjmP8inUnjkaBNer3oMZnxQodOos9LOYE
XRkDDx2eMg5mEXPoMhhq+xVgc8qSsri2btgMAcbOoelaCQP6qSEep3cV6B8VvRz9
Or1NwCO1bRgh9R0KnM+kxzy/wBp5QXwVdTLbSxx4PQsOyPmU2oYZ1qLmEVrr9G4Q
WlCqDeYhkVajzqGkmwWnV6tUE17dbdX6KrFv1n1vaQJ5a38K1PnKXpBCOQmC5hic
xF2VmnMxuC7WtxXHJpRk4slCuvc9HeOAt+VOhV4EImSqEGxDH6OIooM2qaCwKVz6
kFjhCnvTmuNMudoafYq3NmUkL5Ml/ITLW0PPMLqcqL798dWqEkPyeP/XZPB27YwA
p9bZRT2bf/vqw2WZdZ0evOn5mNCN+UvROi6N1G3rjoCrHBCby+xgYWxKJdMZtUY+
9DOyANTiwe3HRh4Xqy42StIuzCuy/9Ohe+IaK5b2yFUwG9kTX9giz+tm5M7Pd3pU
TzGOTbyKthCrgxRYXaM0prgX1xWPeWSiVEs9r2OhNICwRMRPgWIBtfcu6myPVRw9
a2vu5T+RZOdLcUZqat2bmUGHEUa1F3YEbaj3YtSkFKVKD6MVgZ+nSvaFb43J9rje
pCqScSt8tFjA1Hag2VVuZviKiaAC9kPjQxfzBo+9q2QSrhGn/ZRHpSZzHURlj+ds
aGWO3+yH/XO7PJ4FknCssGtT24Em/cIp20rUXzntNZ90abL0miNYZVPYkc6+dHmn
J7vHS6SVAIEWPZJet7546Cwra02OPRO0C0OBgo5yZeD+tq/booKz6oKBNHFKz6E/
sZ/fogBkuuhNllmYCAzlFTRV07D2P3EzBNssDQ2C1FH/E3yDRD0NTnvJAupc/PcM
Iqh2Aai/kQTm8PkvvjYfboZV/lJzZLgjTOSvMW4ENz5j6doANFag/Et4QdH6I2Vn
LqBzb7zCAAvglKbuiY2BK/f4lrGBup/gIumk5gt1KkVUTbe8yWEzSdrNffPvgigE
ZgMhCEx/qUqPmj9/rMIsKb4BRojw164zfgcg+gEmLaK98Tizpuu0QU2d4dRMrbGi
rM6cOTahVBkupITcfg1UmUblwNVVM9xU40Pi0PmkydFAM0I1D9E113s3qzFJO9sE
6rSCwRagIZLjMQ2MBvQWEou6kDNIiXLfwVONlWP/9zgFLyzut+SCUltckeaK1+5f
xbfbc9bKRljRKlfbd0d8lrnbGM+NDWr+qA3eKS7qvR2kEXfTfvoqFDLorl2qGYaY
zekIfDbfIzHWWGa7npE2Fb3gyFM517w1uA0MDNU/8amyHAss9paoSZgyhMtArH/W
O/vPg5TOSep+hGBrCSmi0XflUQ3MFADFNq9gn6Tb5HUv1ahtf/fUJGIJynY39ZrD
4VWHX6JfVMv7xT3u4tjnYQLvkp8iO3xNg5p6bjQ89wgfDZqYR6RsAPhPrDXgLJ3+
GIiaWSpCRvtVY2NMm4BMKTP6W7UPXhtYRAXyxG+hNsVIxMiLd6H8gU5IobfZSPIM
W0QP65pzeGYwf67Qx9hnUrHgI7qSnL2J0VX7uOMWSd/iKaaI4hxn6Gu6WUL/zBlQ
C0q5fuGMtq+QnXteDQCpByGpE70T/ytTQVWAKQsVIp8++PAtidDQgyhVCqb6fHvA
T2TYP2tJ8tvZkeW2apBIhTmI0wKXiP9tm9SNXUXFuIgS8oxm/Ip7+wSQxzzJHl+3
R9vOTyTUJlvB2Z5x8ETGx+/LqWCVSr6kmVkgWBluldZLqwAbpdaS9ckdN4YKPocx
DpqyyzdrnnSGPMXxnlIFeOmOp02vFec8vadS+39uBPAPUL44pWFrhJxbF7R0dBS/
oMH7HB180JgyBFtlOxuclqCJHyiy5qwvsJ6So7rBaKcw9MZJS8NIPuSh/K6LBul2
es28xd/gt4dYW8UELwJl8vFY5OOy9S6S3JYOxb5L08QAj2TdOodhiSSG4jhiDzq0
AEj3mob3giQAKMAf3zI007gZqxC6lz16Z1bsGaJLjXx5pdZqQqS9noqod0YHfuIb
O3rqhuXB3EU1aMhiY4wmpXOB7g07/x6MOMh3F9Y722tX33iiZ+CooJSA4yAcXX60
qIBn5sQN3aLSAy3UUad9JtX0pkhev2/Igf4ZWRKMamUE4hLNujcHX1Y6MzrbirHV
+HldkPSaCPQeogay9rlMkGqvqOrvgbYo+Z+K638MYgiNUDHeyb0AivobEz0CXsCt
JkofnBB/gSVl7H/pk+nuhteuY/i3MMsXBckk0hUlzDmna6bIG6UMgFrdxZdLxi+o
bvlLWu3zBWQBiv2/tXrc0tFlh7NcrVF6weVjrKSWCjwloS5RaW2Y6HXsqFURE2z2
wyQhqt5ZdK5RNktAofGY/RjE21xlSxo42XFFdXLDu5RnOZy0dR+3+/zCxuW8gXos
X1C4jTdVCgpNIHFVSOrT/1e+C9S9PPdhsLRriDGYkEhSnQE5o2OCrSYlRS/srknu
bELkLkQiXkA1yvkD1Wju9+vB6ngkMa6I9uf5FvfrNTEYnj3bm0NgI+QgDIVJ6oMH
a/F1jXlhOLYtaMJsX6RLJvFc2uvaOiNaH+SXD1BkzpURJ1q63KA/Cm53FyMwGCZH
Q5OBiMIWJVCx4Hgc6LT/qB2RKweNPeJluhz3VCzrtkGPF42omqvH6q3Hp9rgm5C6
zZNSDgY/aNYZ5DnMea+7cW1+XxNcafemmVlxP6EF7JLfRM2Zax3iQ+sbGjauqAh2
6t1OEiH67ybx5I+7iGgnins24z2v4bGY948ysIPIG0SU6p4BWMy4USn2f9hXekah
znUT4FdDWHt/3XEW0T+YWbpsX8e1MfjbE1Ap3iRER7uD9ySjJfeIxvy2RhW9HnGG
z/gUCzIfeVIJzRzeRZXxXOTl5tFS48taTd0l6+6e0FJnUme2g8OFIsNekyLSMXi9
SCdrdn4cKlWklZ6klvoBZyJsg2ducUPekHbWDMKtK5iYYGA0yBTBuhKyf9zf68nU
Or54sYwTlEG1/52gg/sUIa8EcnJELd1vNKV/K3Gj5eRBtx7yYtG8ziKzmOO+Iyar
yX7/IBI/7dmlYrCfQ0tSmd1m2Gr5UOmqG3Wqfpv2OT1ZVfJb6qeyMRb0vYG92WUe
A4UwwIcFWJTANEhyT639grkWpKHq0WGvLvPqUA1k+M35GQhFRM0nN/GOXyHOkujQ
Ua92XbQqdqdvSHS/NQos9LTbpVHrmWywQWpqGhYW7wYbM9SOAmeCEAFKF8uKxxxQ
WDsan+88HvJtdzRek52SBhigzJ77Zr69LjJGWHC8eqJiWJnorkmKswNbGqVLcIWF
rdtY2HkeSt+nmpOnKNsXZcN0MElDWl3CjwHHY8XrnydYmEUga7Kf+bOgsRKJKLq6
B5TtXed9suNw4wfj+ZU1NjqDs49xg/ywIgGgUwSy80dQ2wS9zkCEXvVsQ/l7krYw
HyraS8pn9+1FGf1FWC4hAnXhI8cs73Fl+o86IFNGxZIYLKK6ncqkG/7UQImQhwWi
1EQyTW3X4PRugThQOuSDajW4/PvUZeK2eNOEJgqIAuHgCko/QzMdbldnYn+ij2zg
jidWvqsu2O4srkO0trM9AJDIdsfh2t4FVcDp+ltlVflr3flFNNupsmWazySA3fmg
ikX+HlR6ZOfpdq0AtIMpfReqbbUHCGY/5al1+66UDDec7o1y6iEKomCsTWoHIqiV
Xl0kRr0csakxcn+N7N7lSby8Z/c+jh77JaeBP2eh1V/q0KId2oeOtmCyynkKuiqR
CC34z+rddpFZj0OTLfqOHm1p34ftU8PAmlhysL/zKZYiB+AQ1u8nt29uZIvNHrZ1
+NdG22DaIOgR/JOZXy9R6Se3kjVS/ldSdOrGSeABHAHVy01/hQ2vtC+C84QtHEaq
RRg/CQh4VW+H3OeuCLRvz5QeNH5PzyLJEhThs5wQlExFTq3Uf90x7WGy3Jvw6f2u
RntA9OPGPKlw3G6ReBCtvKZg69ouemCSXyIt4N1l3+FGjqnTp4gzsf8IwItZilMy
G+QZm36TzFDvr2x1AXYAHHdFycODIPrhYPt9kbqt3WOY7TqwYA5p23urux68xT8+
huUBQVHAqEOzxslwb2BgMRaxRsiN1eBZRQC6kcbnynNabwxccwaSnMkyRUBuqWo4
2NQLALpMZVq7GDYD8kLQ6RhNeTCiePrY6eCjxos0erLHwBO2kNtmBMIyuE8udZ+9
0mvZOEVpWqY86VTpRDZDllGt2x9qegCh2kxcjNZuKTs5bmjupVlJuxHsGr2BjVJX
7wsaSQi5SpSbc1quTycAwepv8NrgL8vq8RwEg4AbFiNASyDqsOi8uyM+YldMWqzS
kqQ6TBEy8H8AY0+15DmMAUPk2jNjuA+JSJI3ciiuLpGOP4PnVYCT1tQG6BvRuGHu
thPadgXhTGece7b/t+M5TVF4ZWXVKVUI4OeeR3/NAE463QscqMQqB8Bpwv1Pxxzh
nM6iC6XwjZfYjjHZ8ydgCdKzbP9zG9XlgbJiL+aNy/7UWyt5WmAwJ6s7aB5O2k1c
Sbrd3m9BLTgFx86HkQlndRjvjHEDf9RK5LvSyoSdoHlKKhkfZXEEe9FdMDwfGa5/
8Vb2jkwWgA1qeimF4PooVXmxd13RA3o4GfyQaAT+vGU4ZGuz6D8CVPr6OR4DhLXm
11Dzlc3uBH5PigfNDlNKMKbnJRHttz0fUs/OSR6cmXpFmht7LSkZ1iWR5nhVjyAm
EIAjQMLiE29MzirPO/7UOb5M6ApYoMDlCyH0OKbSZlh4t+bGz8NAeHyac3Nm53Nw
Fa1H8JhVOd8bxujQ4RAldiXaVyQqfPNOSDev8GS7+HddeAfBOh+75nZ9yDxhrh3e
LYVrg2Fna7b9nGQ0VIaHIMsObAwGyIfvtbjOwMhUDr1I1s0l6e1Sl1J6/BUaU2/k
OBqJfL38/8OvI1I6BgWIiIjdrfSpRLcQMAP9rS2nCuS3fRr/wU2NOTxMxctseppN
9d25Bu6m2AOHubuKZvytUqRipAMqrBz/R7eQ7NtVbakG0FbgSabt8SxxMgYpWxVa
TMpuZ3FzOtWK3AiiIR2jFHm7mAOYpTSP9xlOdwVk2Uo6SovWCh4ceiPEOJPL4bEf
y3dGx2hV5VCR8wmwC+nXQq+68ivSUiZ9PeETXObhnZG1cXPatdIn8gwzjyz2K/SP
uoyqJUXgmpJ/4zScCRnju3S8Y3QK9qTqRh5+SxhV1GUS8iG2jMWgHEsgTjhksBTP
QToEhsIevzAS0ZlwyT5d8YlHpg6CAJ+7Y5uMAVDObdJyJYZqs9wiTAkDpfWwoqwD
RdOWNAUKkgU1+dRI+dCidtCvhOBLxkBOgtaeIAVBaF3zlHOGbzGx+zDPAcp7Fwc2
kK0VUg78puBQmDNfz9JjkRyMjezJbbkmUqkVnbYF1oWN4elDSfJ75F7PE1mkMlrF
8GD/QB3rzM0XPowBV7AgJfTvSc8fJGnAuYBUzF4B6q/67vwITMvmg/Rhafoj/Gh9
OyOiTYcgPs3Pp2DlBBh1zpG7GAwKparWAujALBN/9y9WRthrZRLVFcXU4MJ/G/EG
2VFrmV3JARXCoYSumYMjwJ+ZDBYHoBW6Op0Jzgv55vhix6bWL2g5co5YqgwFvpde
fPPMiYaJoGMY2vxaGsK61S8PrGe90AJZh+PA4ogyACIv62cPUnfpBjI1JTsukv/q
RJvoBKoasYfYWummFBAgT5nXcqef4Bkjr5XQpnIdHd6sFC2x7QPYiSMoUAOqz7jF
63Ldl9tyu3Rl3uJ6jqU6d/CCKG86ashOcQlVDJ9WJskDqerhKYd4HNiUOoJOKFBn
PpaNqvel5UcAOTCa/JySsoAm3wTW+7e39KliUmiVJ4Ye7bA9zh5IZ46PJz8MwFO4
KLSNy2MLy5iRl5OVUPj25Q2lnJpEwhHAWbqgdAqWnA70DQGsrnChANSxzWpYd73f
MvBHA+gTEJd16NIOSuSo7zekXCn7nX2mI6NNYREMpuPrBPPuWVjFULvDWjj0ngm7
h+aD6TXuI62nbEUerTs62ctZheogcsaKlULI0+C5MHx6LpwxSG/mpH+JWqwq1/7v
2P9yDfaQulqJmQTplbj6fwmHFg60IHNSwh6J5lHKH6OwmK/h+bOmq0esFLcxztbk
uUTLIdzEqA6mbNj4w19G9t/GHlXlbfPgSE5Suhthjr/zUVBgGWSopOpkjV66S4w7
PIA/n+AWYHC44xB9oNzUjRtM+uCW1hZS/zmVw5ZueJFru54clSFx0tcbD0mp+GbE
bo1J4nfcrk2Hpzmf9cFLeW25HrqKJFNigZxM/+Ho096mKS3LEXw8OdUVGsEbuaFg
m5dH7nETg/YBBMY5OEp4FVyjNwEl4hGRRpyyhQOX/VxnMYueCOe4FanVYOp0p07U
/PGD1ptW6YJ38FrrvlsnpSyVnj9iF9cJIct5aoeYbO7G2klyrfWLX6GVbBZ8EQ4i
1jV5WKLDj5zyno2UizGMwHkugWf/PGQlHojpPdpNhH4om8F7C1ZmnR0cfRT2QeOn
n5o0aN+NoRMnSSDY+gc2/EKuwe3FSyKZbVSIA/dH7euHVYATYjNPT9KsFMcPnYk+
f7fMkxAdCpMTR/b0VNwwmoCS6u40OjKfdvqc7sY+qMfqVl7LmZd2zD0YuS5BJkXA
2hDPLvT2jgAsxSvQNo4Jq3CRrrps55JEoHZy+M70S85NNvGmuXDAEoIXg5ZxiV95
dOidmCouJDYtb0du7fOj2tIJrj0WWvGG1N7sojKZPSgMAzBGuGhYVewNDDdGpESs
v18/xB3MHMcChU1S7dXSTQKVsz9hcVYFo5rJM87ZrOrPaHh10eE5mDqTgozmRw02
8/TTsfcaRX3ZI6VrXQhJpU8GN54pAB3cLf3hHWSmoNEMFMucfIR6L4RWeU82xkNs
gZ47qprOEejIYPd2STx5SvQYByN5jK5ndrcCikW3j38mG7Q5wyQILDVeRhyd3yWL
XfWLKGuNQ/lqVAVKmBC7xGOtJq1+6/A0hovGF596Sbx84O5NJz12GtvLowZz+71/
arip/+3lkvAzlf+BjAPLUNRW4ySzJG/S4uas46BgM8JtTVvDUZQo6o4CUsHCRbFB
u9A/74XOc7O67LC2oATcB7/9R1gEOAIrWsJfFbW4FgJAj1LZQBpEUqjtVCsiTl7D
Hz4kVtntfHswiMVP0t4vjft4m85ns+R4WHrazxFb35J7+QDqYFuvDy2GUiMzPN2Q
nPwhYBvgpNs+0mZIiYOLCEetr40x2tCjrpPqIU+a++YeEtUvreRsgYyNW7TTXfte
Gq0cPEa8+Vs4bhJVVIPPCe9ajgexW0cainQjfkClrIYphq9N/hLf/fDvfBFTXwil
QOXKQzFB3CROdtlhje1jMkGjvTHFrFaPCkwBtCLd9rPGuSMDzScuSuHAmz2NFKy+
BMQlSYrIPrqM05yj1m6byrJX/yCnQ7z5fSPwsaYsNkXujv1nY7gdPi3EdOIgkQjg
gUeZRS3GLflrt1oAWm1anGAmvzyxqbftGlPD5gb9gV9bAS5EMpJYS6F829fBW3sb
PnLRv19mbZhELzfV79gzzU09Gl+xhBhNqltOJANsiaWx4PxShmVjiaXVSsbsr16K
NWTbMuQro2WbWZesjwtf1a4yTxymkfB4Rqw4H0MsmIEv1k5acnTVyJ2YO6nIzrSU
fWNziLHbvW8h0wSGqxUutWcu/WLzPa00nMpwmumfJdwmHoJ9hkbWuLRfhEa83rPm
I0KGjN6h0R8/uKs2L6DZkN1tTPoYQS+2vibpVqAxzxNu3yGzc1qMXELsLJZfwPdQ
ZJrJjUhgamVLPLg3TMHXIPF3rP+X6x3iAM/diUHXsPSEkh32yz2+EeUZywY54TDq
iYm11IQa2J1OCs7+2wltnAMeTXrBAKMXdPDk8a4V+8CZRbtCk1uk9e/NHj20vKXu
s8zvawyUuteYzNh6pj0kWOf/N9CgIblgiEPU7xDt0JKSYD8keCO5CYerj10PLvZ+
WlFMxaRGsb5R212XhB2UChDMbEJqsRBJaveKLN0jr5ulzwCtnfMRW8D2nYVyHFxq
2P89CUvfhA80pcsJ7WYWHTVBq/CDqrSdTQNjLHIMotcPktlXxJEFaUoDwKBTvCND
3bxuvjtXUtpznnl2iYTdhSSm7GaqdxQNOP5dKqX7tjjP/EtWVk8TeXq3M/mmxRDZ
NWkcMa8omkdkyWNDqdD+0yNLM2Fuk7ipsq6FD3UElp/nX3n6B+5t+KJRwd+6IwcG
Wrk/jKWayzYKS9QaxZpfeRF2/KV/cR+TComLi/HPhLJNb2g71LjBvLGFnnGPw+2O
/+mGJ0gZIviuLoZsa80A7UgjKUwB3ajAKaaiCohBe8xU5NYzh84zgzM3LP5bvZWL
vluESjol35WxsNjap76lvoqgZ76xQtHC7ancMQBiCzy6QOzJj5s79M2RJK9BkLk8
m6aId1vSJ8wBDoN18oWBC04uPndaxvUp1JhgO66uWHaXB84/BViaNLJ6mhxcbTQZ
PE+xS7hnQlP6FtvSoVAovGFXl8VJ949HXHJRxM12Jl02L7IVFE5DPx01n4FY/DtE
jYKYnZ3rXSPPOvzWdTShj02jfMaFFPX6Qav7KqnePKgl1tz6xPU21kU13ooMgmTc
U2QNb0MoIqb3cjJGlQ3w2sEEsmapNfE7CpG7ZAQ2Igv1HVbxHwIGs2joMkue7hvp
aRyWNQN6zEVNVtyFO69/Sjk17gIsGMkBiM/QTVRK+qYDL1NNDlCSZKZfnxej1+6/
08EefnZZRULVWyi8bQex0uTPXJsbPB0FMgmKcZeqQcFnkPH12A/sWbT7b/90HBRw
yCoifTetQx4NdL/RioksMgcrVsP0nKFHEeuVkKfrGEfeuJxRj2PGiXTqC0sE/CQ2
60rH4Gbfz76DjcJ4Cfz9Upq+RfL3MeGnZvsdJF2soTfF1gyrYh7kjktixckWwmxp
MwPGtnknAlGdLcH6WJe2odLdtuMy2vzGov1e+2K556mFR1B7/SZYhdo0WlxY5C50
WFHn9fi2w4ONiNt5RMBKzYeAys91rZcIsGem9PtVLGYywuEcf8L8xiv3rwjTzrXI
r2bhAUWCOvqO5k/WpE3dtQ==
`pragma protect end_protected
