`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="galaxsim"
`pragma protect encrypt_agent_info="https://www.x-epic.com"
`pragma protect key_keyowner="x-epic"
`pragma protect key_keyname="rsa-key1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
P1YR2GLJ62bpWCp8Rw6NHnV4SvUTGIG3A6ZlTz/YMrr7/wJE6eq7HmKJXZiMqHdb
IDD8d4MJV6Mrw0oW2o58WFxX87JkCnwcXzFDQ4/GQqk/W3+rgqqzLRXEbyr0x6/S
DTAsf2V3L1VrhPCpa/pQEGKIgDOGcuZx/00BjOWewbRybe7sAD0/6Eo5l+ma1NpB
q/ghMS01fATvHxAU0bw85fbj5tokXhepZJj+/W6LwkN8EQDNVvGACzvSHl1E+1mu
uDRRHn57VwOCXHEXlBKcidrVVqlmoOKZG1mTLO3B40Dafb5LZrwQpmVD6kj/HiJr
pldfF7IOfvSaupZt1Ry7HQ==
`pragma protect key_keyowner="Xilinx"
`pragma protect key_keyname="xilinxt_2019_02"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
FKYfNpaJdF7XQ4Els6uFCVVyuBYfEX/8AzQhkHTfjPuN6wtOijus8pwvuLTJVP7I
D1DvU4T57I8zbgrS/QmFNhK7nwIIjnp4TQP1xP8Qi8ohLXPEqObsndaizEalOYI7
+L4w8sJwuNTT07jjABSH2cMwAHDjSjSg/cjGk9f0gQJRtagzxBuiUoYX19dDol1M
Q6S1p9dhztjgnO2ASUIz86yZ1vxShpGPz4iJXer+jzI6XiFjqv1WD48pdqNc2krJ
Jti6EV4tFYAW3llC74rbSBAcxzhVSaxzhUmxeu14KuuVkQGYOluhCUwuni8+cRWG
d2blZkZ8NZXt9Yaayv2Fag==
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`pragma protect key_block
SM5FiGbAwjw4JfLtRkBvFaG9mv+Vc6/VvmXXbmv6uBc4xlrsAmMG7Revsmsra7jy
IM01yo/GDhILfCURyg5f25Iw338fZUa0Ur5/R7hJFSQtHHWhR1hD3HhJjZluNQz7
cvtyo7NaGzHHQs0aq8OAGVkVGBe3qmITR7bRhPd/9hA=
`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
aLF36+z+RDADJ6ltmFFqiTgc6I2vpRpqdg/ZkRKLxWhP6ZTQszalJtWemZ+TC22x
9ADXloRGLM7r6T6ueWV2L294x1aEIF1v+RmNFEV78ezK85lafckgDLMH1kASPAB7
sju73q7SXe9fSsjgvwk8T3a1zCaGz914w/WrzyVEMrvV7mx6qp+A8hpOOsLB5dCg
f9sDdYVB+xLy83gTnlc2FTazNbtPCXOvsMZJKGd+UdNOl5cuScP1ai0+87goOlIc
wNagCwX5ZHxeFeJvJMrw+3aLZ4qy35px16upTnUIDmVmar0yl1q1nq23+PTImRDB
T4WyLMYAIati3ABcN0hV2Q==
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP15_1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
Ayok76zWfiHGQIrCyXI8LONUvuTsRoBemESMWrR3vn2rJamzfDHiuFLNh9afmLED
3KlSK0tLxnhQAE6O4RN5IaC7H6vSIDbcNZknpTWPVTnNOI09avi3L3CV5yY2Tl1L
Nqn/x8olNSr7+pzvbhqGcsONRsehat1FCg6bqx37cAirzWq1Zg2L41CprihGkwPe
rZjiZ/g8+00/unBIx1kc0osGndtrGiO6PiBGJHlSKk5Ch7bQN8/dP6I4oCYaZ0o2
xT2qmoX4c6XdLfjAkpfX8vewLF4HdfxykGR8fJdn5IxAlmZjbDR/9Y4hGttpCIwi
MDWs04xQYEx1MzYkNGsrwQ==

`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 3376)
`pragma protect data_block
KpJ+uXsaGkdk4CD2aUWSAWQLh67uzME2D1/p30RdTRusnGFTO0UVrabJwbMWBfSM
kLNcGQkAsy8Rsh8VN2TzU0YS7KhA5OwOn+02u62a1WcvqEGpe9W+cDsWOftahf40
o1/3sHxz2Kz0XBuqBfzQXCHtehdR/ylVutKRvIzx7rYNaL0/DkC7WgEch4SlA7ua
nOEXK1zAffR18HUCfisC7OpfvA3O/k/M9IJNNLxGMgHRum3K0VPFFatxWfXt1nXN
wi4V9iWklI8EleV3aojNTZIOtTj0RZ5HjoCyEndgGY3XAhJh+PRq3FnK0uAWvFmK
E9541qU4O87YybFoPVH34WbHHlNpSnpPUBVBR0bCieyiK/kq2DK6hg+WZtV5TT0g
PCsUz6kCmL+EpiJJQsd8Oua91DowHa312yabmlSSd62W4ugC48tDm5knXdPw6Li2
2HdFIca3ZAxttyTKjxbDucjKwflxOotjvIoPyDO7osWyFkj64WvI4cnf0ltj2cSD
sfDsaWzFVnb0rirnUpwp6E1/IjAT4Y/PkPCBL1Sv5fGcPv+RzUInNAJCAOcNk6mx
wF6hVcqYUSyUetM+HIwLduriaU5RR30YaqDfjdG8YnEqobznXr8LX0QhaYH2Jfaq
6wCHVbFDage9p41ZI03TRt2XEmeq/90DFSqzVd0qqcJaXjan65noFNRTOXDoEkTA
PbepHQSKGrA4yQXozA+RW5ic7XTiL69/w58QAoxGekK5DtuB0sf0ek+gHQif99yo
7lkzs+g2oMLuoewXz2+G3GM7xrAr1OJBsgwWhG9ST48EILjAgmf8xjDM7Zf3UsKe
4u5GOI8+0F1RT7gHvJuhAGFUN7jw54PUqJm11CmngLl03j2moXgUls59HhuvkNih
KwS+ururUVyiBvab39dxJjc/UGkSBJ+EnCU0hyZUhEEGyKtIssAEHH6GOv75x5S+
ymzdVcsavsHkrQP1ra9yVo1JbxVEcPbaE8RqHK05K8ycmGdTyKd1AJJqKx+WeLIB
YDvuv8xKFbx7CKSzhXPILxJh/plY1W1ZY3YCMco/iDoRoJNQXgAUeblDIXddaKE7
CgOixZdrQax6WFWmeHGFyJKop53GqQPqeUaIQtwAC+MJinwE2/m6p/eNcnB8eAUu
Dvchcgnli1b7sIley4TkN/i8P6nCLjH3k2Vf0Hzjo8/ffSROm3Jq4q3Q4616xWxd
eCkgebYjcVseoCEHaSThgGhJYWZsan3Gv/ixtFvlrE+JuTxFxozsofpmVdqWnVt3
rP3Xpa+Mc57JrVyPx5Zw3DOiv2sj9Ecgskbr08IwV08PpJOh4f129BAeN0KIViEk
T/yhsRiOxAfjhBWsPubdDHY+MIKsERFtwAOKDqQt8XjoQNhRR/y2cGXkCQSOa/hg
JHzH0NUqBO22x9dmYmdXwXnnyIthH7Sk4Hw8WQ8SmsuQcnrcCGb8tz5lqYR4XpIO
auZb2oi6Md402429moHNl1q+uvbDSwj6iU9S9nNXDyLQbFzksKC26ETBHnLUOKXX
73sRUN+Q9vzU85a35ociP+GbFdhtyQILEXPI8XRbQmoZvFZC7qUrYTo7NAHDQvmx
fKZzqHF5EaHs/JrlWWSHOsbKcx5p1XfzL7Rte/KAJpBvS9PNwmaSpFEPKtUHEMth
MnJV1HTvF5hvwfn53y0MpuepcMXfVKXa4qtM99oJWBKPvIijEsxrWJp6mzRGIFfi
EjeszZo4qP3QSzl+v4zZJ3CAvV+1n2hKbGxNPICatL3ol43ANnD3c5vdSOwg5Tk9
M2KvvjKbtKyVHLRXi6zl8St6tW1aU2CklkJ6W6Qeb54DmjPTbEMUn9sY5pt5Tn5b
J3rijPeVTip7ZCiFIuCqEM6wdSNjeOAyBxFNqJCuEwyXMMe2LuPGuuiBXs3L40b8
BHprgHax2bdGjVGlltlSQu+H0CcCQl98LY7CDiu8znpIOLLwTMb6Pf0i8RU8dEQu
V00BjReHbOe7e3Rv4mrhn+gSeHxQS8B7Q9X4nSAnIQyRWh4Tpa0jBTNsL/fm91/E
vA07jUIKfxgOpQcLYkNy1Ba5nUV6w2lEVxaxtkbE+rbZTqntbF7C1KUG3IigDF57
I2yaw4O0+BC5KSM1hG30dorsRdCy/qfFT6Xvw1UTiz3R0BrTXb60nznqqDUwt04c
F5SV/pj8yN8F0dL9Jzgf0a0IpwS3Tl04SgtBu0j/iRLCjhBlTmwQxTbr/g/Wo8Nr
LYYvT3fwqfAc6TF/QzbwXn7AqqQ2d2UScibaWZJ4+f5NgazfjWCD35EzswPuD6mE
aLnzI31srTihsRn1e5Bh6tw6gNLjEMCx2iHJxTme4+it4LVlBL5RbksIPcf7if4y
xI7vkAVHPjzMdkr0rBMzhrIriq0qGFLC2v9dWoxFMixuJeT02/XTSOS2JdHJgevH
YdIc47s+nclAX7XUTlVsKE781a2dbjue7TGomfnHUfb8WBkD6h+/ca+Z08CJ2YjR
fOid0CPEBVNx++jHcOWfglgjnVq9nv74P4TdL8lX8SnCG1D4WyiJ0ZU5GZHzw/Uv
QXHwxQczvw19p0aW2+xJah0avs3dup0L5o/+kqbqrCI0QIXT6b9ChsJ2UkPbU85N
QI8Dl2ScC9q6dQk6Ggb+VzU8VWvd/pUrfc12AuyiMhiRZZgOx0Iqyht28hzRdCwg
MlqJGdaclGIpZkMYng97euBWvZGGnG5dwzc2A/LumBEHJ9vCaC6M9YzS140guULj
PA0dcst6/nYp4vlRFclDxC4FfLFTiMeD9BmKh7hH+hvcjb1Jpgy1FDammlfyXyYK
WjQ/Dj+F+DKyg7HI+qsQSX3wLynl5GDkaxt6/4cRKlOGoSWiypKqDidiLrVgl3nA
zWJWXOLhTahA0KWT4H0NxhuBAv8Ih3U+Jd8Bdof9YHALUQZsGp0+GiOwB2qBpHl6
xfFQgkbs8pzco1DNPRwpdgRZGcgZDSLjf5AIeDiLrv+nFPusQJ8cdQWsM2GVXxj2
lh/CmcecFIpR0Wdd1LVMPubrsjG/l5j4eSpWhJYLMcgFMs4op1rM2C3u+chrAmY5
5/LG9lf4hzpiOwBV+rIMb9aEPfjmacTACjadQkYP0ZjJ5MWYBqfFdQAaX/H5Ie+w
+6fQweQ83oYsa1GmQbNFW6J+4LmYV8HC9uHY9SYbs9N/jKGpymss8IMujDHQ7gJi
rvh73NlDxTvaG9Cv4t+U+nP1mNLTdRHnqPGEDQ9sZQfC/5jIU0JwwOr5lW4+nbGc
/kkGPMMJ0PUVHqruGt2NR0/dm98UcmAGLiQqumIQvAeIGifWqidEJj8fOTGg6Nzg
dXLUJJjtZaViIbwr1IhuMy7PQ2tAMkgIyE4tYwkKd8B1WVEMOKzrs7mY6hIp7Hk9
RxDWYfST+6+hJvuHp6bqqREc3t2ukdNEzL5TICxM51EbVYq7x3aNwi18y40lFYfi
/lebCET8B2cvSMi/cYQhi8RPkmfL7H43FqIEnCcl/J46BR7khwejRPyp1PNYg0Lm
L+4xpi5wDpky8v/piVGtGrxj8NKR9zgZFlldz67xbk4sveA0BudogGOiS8eeTrJi
V8EBYZ1bQ5JdiJ3YjDZsYZd+qlIAncF7QECQz77vM+LgfUGrkWtny9g0z+yA/Sf3
Kwmf4CEWbhdJtFUvVtZz6EFD09Tw01m5M4eJgXBD0N8YHTPsECnuUxIH6e0H1JMZ
BAXjs4i8fUmEd/Xpu9J4eMsXsnvJQiaMY1M2jDn3/ecNrVVZROZ6rqJrMOKrjJDU
rxOrfg1ySCLvpiAxeEkkDHkt4huE0ZyTaTntDnGEfktCrfGM4sNb+8SvT8Et4a7D
8ramyZY8DXSEfoQULBMTjqGvU4qYu4a22ExTS2G9KgdmdpVXTpM+v65eQE3odFiG
TBORIJTUI7eXRiUdtHybNi5UX/vwAqREXK3jLWkJfSe23u+AxP9dBkHguITYGdAa
Dh+XxzNbE0SoN+/zOirPY0ghgHu91CNtXKDrFFNBn6jXiFBI/bc3uZgvcrszBpWU
PBAU+Mt+Q7SAVMTjnm2uTpIEgvvE75Va7CcW2lo7+ynxbAemR6InW//UQduJG3XH
lEx55B96ggwocuCCJl2W/ksC9RnpaAvfMhFB4UB79e3SyaOVgJBrKuSv/LSFLbCE
eBrlOdure2ngFqpAQCEbPE6/bjg3DYIqWTZW1uz64P4y/j/S91b+5kRJQ7QVxJ96
AGwLqOVJvxxoeqxSZ18WTlAu5IY7n22rWPsGCV56+wY9F+MwSeMfzgVizpLhJjiq
YufhrkIGnV/IT2Nu5JexnqZRm2XWn/2U4MYqNDJbI88qJ/H+5w7wBmkzZeOtGkec
oHtUH7CRgYZt443XKPRsL1zAZvNExhP5oOEjVil813qSrdIL3Gzw7nrS04EgR0xL
N6REC1L2jeHwswm11k5jn3ldsM8TNyhBMW/JpAi/iD6e9nfbjwlLraRR2AAOHihD
99hXMTEq3fCVh7cTmKF/eQ==
`pragma protect end_protected
`include "xaxi4_slave_emb_func.sv" 
`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="galaxsim"
`pragma protect encrypt_agent_info="https://www.x-epic.com"
`pragma protect key_keyowner="x-epic"
`pragma protect key_keyname="rsa-key1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
KJctPtj+9nlzwL23dbiWOG5gI5yaPEiY3CdZ13+5B02HRJoiitUAAzMsbkiIOs0c
wVB2V+weFG2vuOiwQgfKxXuKxPLcO+dN8hpedNCYbWkxFi7anIB7ZjKdv1ZpPOXh
O0SNaRwtp4QoDw85Wsr1JNDNdO8psVzWsCvNInF9yOD0hNlKkIt1uZLs12D6Uf7f
WIYiIYRc5eGACY+T4eCnbF70sBm034xAb1lELxUTeWSwaILrabrHgGJSDPwTWEnJ
dPL50jgYYjsUnNfENErl7IW88DDQNXQFhOUgH5wmyu6Cdt35xlw/HAAVPrH9Byhy
+LWvh6DMLkZ67GBd2R/n8A==
`pragma protect key_keyowner="Xilinx"
`pragma protect key_keyname="xilinxt_2019_02"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
RP5PHB786fSZCshUjMHguLe9X9iECuxpiAjbsEesPsmUVmbqEP7hVwsf9yi1ALL3
n8UUIhNVayJxEPWxwuhGGFQNyUV2vYrbrLumPf+Da9XV2PMKuEnognpS7EVmgEhV
xnu8PgvYct5whotbdiOpZ0qRe9XV8pud/o7rBaabZmIHfXZpZQtA3r6koM3cDlrp
8B6SZrl7RysMBESVwxSHAtzDUcSXFuWwFEhlOM7hIezFSTKIvhKvSw58jPpsxxGr
lTvPk03/nO8XkCGPSO4WD4FkLRXUtqR2HB5Jiw5tB6aaBInsfYhBMkbbPfZcW/aO
EjeNM0ppmBtTZADxASINpA==
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`pragma protect key_block
HILOJ54qPs25gMTGZSQZWUWYBSupUihSSpaY2W3EYXuWHvA4zXNavQ9Dr8hahiLV
v/aB4FDFvUR5M5xh5cdBkxTM6IuzgMunWCb1val8HcYM0IhGYiQxvbnK1SdSmNDc
kyHmdB0RFrlfRKqvDP1nxd+ebiwbZPJrKGxcfMnrSJ8=
`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
nqZ8l4zlNJgYF2Fi0Bz+UkA68yNkgPbMosnBAMV+acPMTMcrRnJ8yJJt45MpI1kC
uaKwVoHBEXbiKsvKAw6xxdu7A0keiW8ubcKTNg/3PEQP0tQxquwfNafhxqJYzPyV
qXX939tgStFc55xMCw14cmHdo6XEJvmnL8n2xLOTFCNDiKY1tbsXUr5iwZktOa49
RsWf/ytD+0ZhuX/pH/9EpmRLtRT804Sfu1YClDVN1zfL7bbKnygpSSorAn4+huUQ
aJugMMfZk86bi+fPBMFPt4PFCAQoH6CyzXWSTcti4U0N7J7wNFJnmYwyApbE4Pf2
1clff2Gua68piyC24/eLUw==
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP15_1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
37wD/5C9h1jqI6mjzRy2dBRTJDj2OuJyqfl+LoSHlaFkEq/qbIAqkNQ9yIr0Xkla
muLh/5r/c74nwPzZy17pO8h2L1+0oa/nOO0TQmp3UCfT+qytYPedq+rbAcX0xgfp
SsBrP+IOT+R0ZzmL+CJsjbDxm8ZR9yvmFYlwILOgqgXEHGVIUV+U89Z05LLNPRWW
SbbO/I0PazH7l1JaV+h+BcTBxIBcIHxpFzpRTjyOxg3O33J+zMjv7K7txk10+jV8
eghQjChLTGEHupWm7fITmHgELfwtbZq0wq+UPwKWs1l0Q+tgbTciBYcRgqUoHJQm
Wh4Cg2tW16eH4ufUYQvZDw==

`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 4064)
`pragma protect data_block
fm+53kgArdglkCHhXULB/g3fqb8T7zECb8drtJLyeQrXcf59t+x4Vnt4ZXqDjgiQ
hQgtIfnkw1OIdGkmKvw8HB45lYBV+QAHq33I1A5LYzuOUo7SkEwA8KtdJGX93TNR
6E3QltYdnp3XEvABkaduU/fLvEE7/F58/I7eWpCrmuKdk3/pQEXp51Yt1al5qW9m
2DqG9mVyp25jpkgp9NoCzvCLVLiltIuhCxfXwHr3DU0MiQRyaZowlwb/sFB+Uh7v
sPnvIrwDWamgNBeoFkF7Y9rbHEdWCgXkwxa+3lANXYf+330DMesb2jJWu1diDd8E
VeqXFXoyuvh3oMSVg4yrz/2QZA9vKb7/uHrNPGkOlyAt+haVv+kxwpWdHX7mlKTH
mu1hBwN8VelUwyZTl/vJiTip0JoJiMu+FMvvisl/xqjASr3VfJrh7BhhEXo5ZSh5
YkzNbQ6INQ/oEUuQ0+9wWaw/RbXb8IunnfTX2reP7ArY45qiYpNEf+MD+iPAwe/u
/rdaTV20M3k6vGyT390cfwOg7tE16nqG//g4MAh8KY/iSk4dQ21yfq0p4WCeav55
RTt9CUT1clqqhnzTV9Nm3GJp579mU5JvvoPD2PBXbnNJooXQHXpAlL7gAx7SuPu+
wziKVmwD7noFAAxYvRXMkljnJ+sKpifOa+++NYuLOchGYAV0NAe4C9oBqL6rJQL5
oeQSH5d1kjWjSCp+ndi1ZFSkZoo5gXqFuFMqCqVG/C7hgvVbJuE/8+JD8Q8jzoBJ
MPGBJHvHFtjQQ6bfobhBuiaqrZoS3EOmWtsXM99+5ZGCB0+0EB4MU834QtZc3Q5a
vf5k9znHdT1E64c7cIgIasmUli5iWVHZU7JLCbR9usy5y23xKDVYmCfuYsfdeaJu
CiQxtviRrf1LF6YjdCLB+XKFwNq1AJEu4ocb9YZsnse2EGOfkEdN1KVD1JxAixot
zBeXflQZEOa8gP9xQjHSv4QyShNGILqNLGdUh/ZddtWDiFEHeTOtBJPmUfoJiOph
q8FwVRBEb2Ps4G9TUHg2r5ATIbsskCtIHsMQX8KaZUjt+8g417UIMIcsgE+58PGR
Ele8iDgFGN/q0rZVdBzKeIEpRaH/7nxN2gR4rjgHbBNzuAqK1OkwNqXhW/T5MiT6
z/RsRh8iMGbIah98Vddws5zWPpP6NC/i5JzmDw/m/+8C3xpP7mAesmO0FBJVMHvT
Jc37hZNDhgDtY32WXf3GyxGrn0lFQ2gqTkk3T6G8ms2XbbHD/HJjx48xrJ/PTTzD
/f2R/cI+/cdJDOZTbdUpE++GvHG5Sam9fBFOwCmo5m9E8scVMFquwPcq6agEJm3V
S1+hPXNsu/IogIWs7Gif4ueDD4FVk/wIRkm6ahg4AeLErpfmNzJj4zpFr9pqmO48
KzlHT07gJ8gq+oVDbSZjurqPQIpvNEXwf3cH0ekdGYVUJ8owRA5bXaXnmA3pDpxx
z3CHCh1pXzLsE+EHq/dDzoK/ZsidiHgeLODw8BI9i7cvixejs3+ZXJWDYhMVeBMw
pG5R5wgCRDhh+GuFMYHyHHZogDorqyrPmWkagu97msdD1VNagO6RWbiwxBCVLRX+
iZ1iHS3l1bgBa2/O58fLpX/kk5z6j0gMPx6EHLWniRzBBcgyt7pVMsR58NkpzLjz
LKIANDjTqZS32dzUzSOLGDRVm0Hzs60lNQ010rIb+mDQ1nDMHg5MuJ5isd8XiZYr
TUbmADzT+ldC2JPL0Xc1vZG/E2OOnHDbLeQJl4cKg3vGjT6p9KUHGqM9ggUEFch4
chvxcpaZAOB36kvGAreY0Fl098WefQ/jzc/rNpHoj86hnUav+Ek+VjcS//qNWzEM
P/6DFnXO0Cg9OAtuLs0ZMnZOWLv69EqtffT2Gzcos5nOrXiwUmI5kQeae/QM+0wU
39p6PoXxVJW5EYc7CZg2O6xYetztd3J1bAbus5lNcKYzVrR5CPfnkNzsGnY+i8jF
0d0qocM7hNwILutqSU8tTM5FQxkKmkEK7qCK2eJ1uvUfVEsj8tmshQl76/2beu8m
M4aQjcRnc6bpe/7j4rnyvy3TJ4Si9yIk5HudD9bESva7Fg/9ee509fj8RoXCDIFS
HYSL0iG9cbQGaijW+peW4dTPltXdDZ8MmMkraJkAVAujvDt+IzXj/fTid8jUuosA
oxzXa9dqCma5Dlh3I6rOjDusO18U+WTs+J+pL4jC2fBa3CyI+ZLpCn1zMLhggUcR
w4DLBtfyDKJq07qrW2lrG4e1l66EcvjrC78A9bDxOW0oLwkxGw8CYz50gw3rMCNp
1n4GunvylRDb8xyLunMIiEhoeALqzhPnb/D3SSfJh4PG4Epto++a3eV2RZmKgZa1
T0xCeMHXnY3gdTlcwribccIoStIBQSYa7GTaH75KXLZOfQ9Cp0C69zhf9XVi37CX
rqT9Q9JSvYJlK7BKFkVgcz3NnMwQ9e2fh6AMgphl6WKfJI8uUwDNCHE/EmSUWs2H
zSs4M8EY7E8prAHh1gwZyMJjfG3frkTeeMnHHq48McKgAy2vuLrIhSyUZgOZ3UHj
ix7s4n2lBkKvxWkT4LWcVim2YL5EqmAJxWcgApWsrDJuoxJZY7pV8UrTNixn9WLE
D5a/DE1pw2hL8L8cHBTjI20Vzhq3mCdjJy1L0DgTcFhTu58bebSQ2+MiOpvKr3zh
WTYKiQHgN40zT37c+1k5VOn62uRHVHCW0mwW/BeunEv9ndJtIKB2KGT72vPjd7qL
4lFQ1vJubhJ+bJGW0N9kcPMTo2SliU9nldxDQY+Z4uzYiqyQMevdanVB3j89z/BF
Ht8e8W8idg51NfUBRvAEU95WHgkYNzUFBvLb4B7DY77gDKjtTq/2LLaspybNnujq
3/LJhcjkuyUu/N4F20qIa8jXifRC+bpqgpuGw59qQWkKpKmuXiBO5rBu/caDchgk
tEVfdZ2SrNcFE1+JQ+CXu4WhHRx5XeC7yCvRjwApLFhk+YTWS8LTcnsaCM7DkzBh
opoi61RDFQ79TllMirLcCLeLjmQu0aO+gHicIhZ9BUlOCOgm124nWO59ffZWbAnn
w6xCUWs48HRsPyEOSI9Tq3Tth2uMkSIPPmLlv3En7XcXs2YZttEemg49G3nQ93AF
tNeJC6G81pJi910xPqWv6cVUr0PKpAMGplSJ6W0yIUxzs46+ZDN6/n9HQ+dZKDbp
CLPgiCIxBmZy9LHyxy/sTBJRVXTRvFKgA0PvhIteuml5SW/OdmXkR+8NELWTZzzb
1awBHJh8Tj5MvSxmh5QIWidBj4dPKh2F4x6f7s3qqueDmfSVt7ctErZT3Zozj5Yd
ztqtupBCBlaQEMmxdcfhxRaVRFPThfvqD1cRQilseutvouNUPQJejQUOIJCx7lK0
YF/W4D6p7KXOtlTXaIYG2x96YzrF/Rk8s4grBCxBiY8VNPpphJ4/pDCga0oKPcfG
1QN3/z+PevBIW5ZobLJkBkUrxuZ3wZtAerRDUifQqQCtcAw42hdQokVONxkzsqc4
w+gYN4QZKO1yt58p/E5nI60eXan83McDUqfCiu90qWvn/Ax5SopTV6OgimRHldrw
DSyMh9vxioOwKGHkPkFwYXtbxl4h/z8wxrJLjZvIJ/iaG3DTuD926FFumipL0m98
mtPCAwTaCTfN03tL8KhSIJcE17U9U/SwUirgxC5v+H9Z3Br057Q8fURpigSREXL/
mnnBltghG5l/ZikFzC4Ymh34AVEQWL8UP+VW7hhMTBv0fRLfG9HGeDyqabG0Lue9
tsuAXfn9FHmU4fkVqGimWb4Dc9vq6Kz7STFpsDAAY549shRHV8zpzQoxybmALqAC
NxnZm+j0OrjyqgzKFAuKZ+/QuqcACaVVDtfBU6kGO/djc+hi4uXeP0d8qU6xW2KC
9j8iBGUZjXQXhFZEDqHLKf7JbQ+Xrs1dK6ikrDt0nxfTz2sDsE4PwKekRJZeF4o0
+ftCG3OeAy1d15qm837cFx80rysYSYbG7Vcjr+Bi4kDnRK5n8LZZifQMOsa11nXy
1Ttxbi7fjWlxVhuZyI8+sA+X0UeQIhVT3wE+6g7ynnL7deHASYsmWoIi1+rs2COm
+uZOmk4Wd/D+JbisEYZXON3RLGGmP3hmivwNdxbLVPKo398kTINLdCcKBYIfqA8g
xUA3s6ulzDhSyiA0VyCyly1ixvEyI1jLn4/c4e1mpgHLynlEdZMuh+o4p+kZZIJs
uoYxZJnocdgRSQCv4DBZWufVxC2iop4/IyoOtoO+2/GawMK4zay/J7C0jtuBwV7d
/A7xGh4Hti/gcassdy3PNORWwLcq+sxcaJ6LMYiWY2nbIhwTGq0kZvE2gNXPXu+F
uGg+xZzgBIgsrBWqWnmZplRCAxSaNihqmNMguZ81ttKF7d334B5T6hhjlGugpvlh
em/tDJfDMY/Jhnl6HmrAtw1EOBk4C4jyyItO3QoHwgQaum1j+JVOSvtp/6y/sh+a
S3o3w8jjRjM7yMpjIQaaOq/Rj4+SIRXjw4JFEsjv5pinJeEbrtNBW6mmSpe3jrlz
6ZiVfAqnLjKGgMaBfX0DgLmdAmoM46HpeMqqxmRONwN48kGTi25pAt1j54NC3dIA
r7yqy5OMXpoXGuyOaImSr0AdDpMgIR+1IfRHSiLxNGBfA64tGXJOXVcF3fHAEEbh
2lRCBk7HlOQkrRDtsbb7B5JG3pAzT5pNaGTr6Lx1F7Pi7oVTjuUn35Wemx/6izF3
S4AKbJ6cG9ISnAk0rai0wdryPkc68QAUUAY9QJD/0e7FwMlFxRUg53ssmdkPoIIs
lzHV7DV9YMEzuEOfB6T7EtH3c66B3UgDf7YhZTlK9Nnd8Gee5hXxIlOQXDH75eKr
WOb7oMUO0rIlGkYbKfEoxLARHG7jndECYi7FKiDtRVeA6ndRxZs5oLQoQv1upQGt
EUl7Iy1uE708Bn3d4Zz5uOzzQraEi9DaXa4Iz6bigvffs0CuuNd/mrsdHn2wP91K
TZjhj8ow45s3zgkbKXFfBLxlkBhWgSW1SbnJq+Dzbv5Bc8HX0pafgy3ljUH9pxwy
1IAOLsZ+kgUmzbXfMBHxDZi22HMlVbZMh8mMoY8sX2zEN5vI2S4WD0vkguRIn7DR
4UZPvyOYcbN1S94t7lW9dF+8x6MBhXuax6otB38jj//stpeSOKsRLlcB0BfsNbvJ
utXwrY30RmotNZp5uGVQwQk4niI+GnjfBG1ClLQPATw2/F3xIk46O5uU1Fu+eJPM
jFC7kQW37OVVV9gLEp50hfH/bxtRsqv5PEUr2jgynNxdUrF8TIqXFx8sNEbp/6Bd
SCj3aPpvQh+GdBnfovJu6GK3degKsn1qxcIJRHKPxZp5j0TOqPaIHi5lxU+fpVXS
ABKIecft6KEdHAcLNhAW36Y4hfSY5qLPVoaYwmsd0z8=
`pragma protect end_protected
