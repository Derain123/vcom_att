`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="galaxsim"
`pragma protect encrypt_agent_info="https://www.x-epic.com"
`pragma protect key_keyowner="x-epic"
`pragma protect key_keyname="rsa-key1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
O/gp0flc7LtWKo0tG9LsyS7nrxdQt2ScmFaLNqAS3VDPf2i+hyEgyCgG4x4RAIvE
I9HKaYi2zcp/tbem3HWcJAY3MGr8urY2zM1Le+T/lBwx0wFb6v9YzEIriWmWKWh9
XGgQTGbzDo0gKq+4O1PSdQCUwNDvPN3SFSSHnL56x836U4iGm0gnYmzO3IBK3AxJ
Vk0135d7jefPUygm1bq2Buluu2wVAufi/RnLPo0zYtMskIBXwEe557SuYIXrfSwM
jYMOF2vUaZ958a6GUjwDhksrnkEr9BigXEfIajxCo7U9U1+J2acDULN7yukn3OOU
cqEQN6GTqHqiFQpvYXHWoA==
`pragma protect key_keyowner="Xilinx"
`pragma protect key_keyname="xilinxt_2019_02"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
AA12LhIlvQZHjmlhEHpjSVVwXCtWHpSBA0txA3slKo2kw5isIYfk1LLzm+vfjvZr
c9nWweEjOsGEcolg4mOAC7ZgG266PQXVOuQtt+iPiSnr92tuL6O6m/qn9A6Ad+3E
KUKmR7gvECbp2UWinvYyq6RxHZJi1KpgYajyu+9oEDhKNo+l1tuwJ+QZEBJ4pnki
aM1KzD0V+PmvVPlcfPjvkZ9dFhGPBGh1NIF48KHBAn5bhRIcRNNrp6MkdfI+B5Kn
jWcFY3rKsMDYVW9D9WPu3cik7P+QvyzsigWmxy9NTjslYNxt2i1F5cwPxtCb1dev
XdA9DxpL1Zj4fiHTjPNHhg==
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`pragma protect key_block
O64k4voSUDcjDN9zx2BiflJVPkJcFwinrDYjDhyh3B5QuYvQ+tM7r2bCu3tFJQbY
I5L+XuUpfeBQLS36fuNu+4sgLJHPvXDzuqVd8eU/K6UkPFfcKmq3SVBsGAlXhPjN
/mOT3nZ84qAE9HaYVo4ECVPz2OuR0OQQS/ZqP3GI5CY=
`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
mfx+MjMzD+vIaVdoDHXVehDYFtBzL6bCFeGcdyi89CpPn1z+a134SEnMqWVEhqRA
Ld02Cm/tF9a1rCes8P+c36oObva24qPBuODYfPwpLKHMkymVtsHkMIRdoXE/XScl
LO6Sh8d/7LcGS7dam/31NXb9qwiP+Ln64eAIosoUpXoVFNIq5GpUIn5UlVuBW+L3
LH0TOgVXzzkAUQy5+G3ye3ENBuN1ZhQBVysfHzTQzh16Vr3h+WKTapMzF2reECjV
sgsTBw8hgg1pbOSwdTaU7KaZjUip2fT0hT7Dan2sbGkMmwUfYfY7U0urJ07hdJEc
kzJPfnWbTGNPZ0flEJ6zRw==
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP15_1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
W3Yov1Vd37ToPgHB2GePHSrk5GNUgb6qaW5ENw+rHQCJdwu2PwRWCGVU3al6RCgR
LPO6VagfucHhOwn8Qe35d26RhguMK4hjHaDLpLbR5poM3xM3VFhCntYVVp7cbB74
crPOMBWZr21ur+ruAILyeBBST0fSZox2oFxh+b1ZMqSy8qjjBL+KoUznJo4OP3vA
MVfuJawvbg6NFzZXMNxwbZv5sfT0Qt/azx7IAAj4CSMb05H0wlFnOijFNR9SvitL
/9Xfiakgxph/fBeHv7CLXF4X9x4QM9S2e/TWUaRFswcSt+6i5S+JIt/z8/IftpwT
NFAkqs5x11tJNEtMCOEZfQ==

`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 1424)
`pragma protect data_block
xMk7xYOnfxmEg7bVKOLPurOEna9SKDak4gapZv+cbDYEgKvB7tfBjzm6neiMOqIp
H0/rPNw85dfxkUYpOYe2PB4z/YtuCj1Ljl1TWeLZD8F8x90MqnKZnmrfFLyRYrrm
7IN9W4qbSXk+TUrjPNyVumyob7fDOJ7pQmjPikfyc8km2oFakF6U6nlGdChBvHnC
hrnD5A3Cl6Ta/j04Ajb+lMT6ShMYoMwW/MpjBn3yPmRT8w5FabE3/PxjrOj+V5+q
O4szPbBtlZ1ZzJ0/N3ZtV25A9NwVdMwYuYfUGD6EzXC4iawe9pzkrWavVfM/LHgz
3Q2jHM4InjkvC4Q+2nVCKn20tltn4Cy66/BU6LMtg+ajadras7OBOXU5wWG/1K8l
sN1cfuwRvS1Jdg83w0Jl8VHkhNyrRlax7pG2TcE3pQ3mtcNzfJjCETN6vb3qS4fb
XbRvJbmeiv9R2osvQaCdsUlyBOG9C4DE2UzyMwlkEobaTKFBCldjw62wHicYil6w
90CN4kctvy6vXxEXNnGfzQvqhevmtqDxD1ShkQQnhNO7woIvGZNSYLBNiAptdv2g
ayAN/SkZ9QQl05/ab8LVjW5ltGl3+YbU8B6bun+IVMTC+BK5Wc3lpyamdFt54DEw
fjJpzl/Zu8JzoQgm1lejhYg7WSlMfU3fGB+yjJEsOMqKGMZN947hiz87e3U8Iela
S6ZsAFYiphKdSheu2mZ0Nf46S6/7b9SkSIQ/yOrFl5DgG/hfZiWkCnUWfBjyFZSX
fiCRIq/6ytEEmpT+ePBOV7O87SRrTI568eUEwJuXoB/H8bCEViQm7wkl4lumGxyb
uNmACG1WfUZKS7o4Z+ZCheoFUB0SRXJVEQ29ygAAQ8bmnH8/xqxVUK0vhhONb2lZ
lAbnjVK3wqKChNLse7Q/uj++QZQuWRaICrpLmKWym31Ogu+ogbGlc2+ssD4+EPY6
+roYKBnwV6Vkxefy5uhCg0V9+FXD2/Sgzz5l4/lkakWYy60V3vA4PyBmFeGT6uqY
BTieuzfkFPVpH2xlQTUVxvHfJft9p8cZVJvApmpXWJU52+jpeR09mozxnMxPJ3lV
26Kilzym9wRLk51+uYflqMVVQUhAtFBZwqCt4l5nERf9sexmWzk/kvB4kW256Zm7
G4oNPBZG8UpYH9TzAczm1u8Wg7XB0Uj8WnMmSxZaXswVnzE30VsTVSTPFqyr5dN2
VmqR08utNBcOPx7c9gKvkUuMFZiw19ulzaznbwoo2cdYuglPVRq/TGHzEs057YPC
5u+qDjtpv8qFPKvwgYaD9+av36E8uJzQzrrHzAwpqiNkQqSb33TDcPSy3dwI5fm7
YgmtRbWbC8HmTeBVMvKOzse02X+rYT4nP/iqMj40djkgef0WUdZqky4IbD+OZ2jm
6844e8GSoud4EnVu5P3ADPv+jKqWgTCo/G3tCfTBKAtezgXTiDBnV/cZvmserD9T
mVPAZ2zcxbej92SmSHmXzFmqSJRj1dq09/gr9B+yyOAU/S9C07rhJ1Ago8rua3Wg
nV0aPlRQQv6wvazw295YZc8skxAjcBnIM7/OviL1npVNH4ZPFm/wZJ95SQTCY/FI
njOLkeV2LmlEVh2+2HoBksimX55eznEIlYtRDkdpcPpg/k7aDG11E5eeWadQkl03
Wiqif+/PQw+NexjY2crSP3FGpzpAMhUzAboRIE1bS+ZiJBI0RddV4eO5w1A9AsiF
FMTsGjyF4stpB61Gu7difOmbYaTuBm6yXtx3YjH/WI3U1eG1uOEiss/islmhog+d
r1w1cvvkG9zIJXLzoxJimuLQBuR2vPHKPCjtCEBd1cLsqz+Rwftb76tO88jVdQjM
74iZUtAfzkk/ert1eFIecUd9GxYf5WHYXMt18xM/KXg=
`pragma protect end_protected
