`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="galaxsim"
`pragma protect encrypt_agent_info="https://www.x-epic.com"
`pragma protect key_keyowner="x-epic"
`pragma protect key_keyname="rsa-key1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
veeUGfZ2j6h2Tnnua6h5uO+88cVcqAnVtLgChlAP+CRBSWxFip+r0uZwQL1JGla5
HwZ9vmy9TQeC6jnJF1gFU+MtJFRju1qWYyBTT+QYJexRzwYXK38ex58vulkciQHL
c1W2mR05DJKeL6HwDM1QLecCA5NM/CTsXxhx9VJrPiKwJq+68Vvh16dIYyWSEWA7
UB8zGrA6KhvbTC8TXmn3GHOi26nGdAiwbHxm4mN8e1sSOQ7pwnRqnomKwgqBW467
lNstAWJnHltdZD0F1efcHBrMFkTLvC/XW4q2j+YI3HLl3zU056fLfWENfIaQVL/0
bLEeqWCgpJvnnG2T+AxhRA==
`pragma protect key_keyowner="Xilinx"
`pragma protect key_keyname="xilinxt_2019_02"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
CW6Zw9mjl3g8RIFRD+gjB5DMIpHTImjqbc+zoj3dW5CkWEEEW3jNknbt5LwJz0qW
xvNDDA93pSOqC6gh7IIX3VIzTDA/SuAj5IV0ScenALPIZ5zb8/7DYpCSZmfh7VLJ
5y7w2UVp2Q6XMKDFSkEUlH0/nKNOvAiSPJ1QFxmgoIbZgpdwoFLUsP5wBwmjMGBb
9jM3AsZl40D4I+U+KsJk0dqKHPGCnrNay5DdlUbbF7VWx7QNWXHSOWCPBTNMhaUU
0ZipM7t4PNuM2HR+nomvpVycX7b8iqAcYzXdkqbEW60yQIwuctye4/nLgU+JIaR1
UPt9w3u+six7UFo+G7BSeA==
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`pragma protect key_block
KuCbtCGRheSs3JEDW6oKHU7DQkFrvrQXZaRCQ/HYiTEqqvx5FeFlt+6niY/GID53
CCNXQnH7ajSc+PxzhAx9NPvvCI6JfzBY8Qctkls3xAjN0eCrGM7Qwm2SKofeLPYV
QBUj7FlIFp99HmW36XxVWHZqothuWpA/N3X4rZj93rQ=
`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
OyZ8lO16Qe7pZwq9j5m9QZPLNSq0FP16U4U2AXEHM7dBp8Wx84KLjowoLfrDIRvL
Bwp9w3QR9aVXOyDvqf+VI/QzYhHnFo6fZ43ESrfnZaiIQDq5QON8DxG2qWV4/2Sh
ErAecA00otya/lfh6b98aYra30UHyatwLh2em8zr5vGMsV9L9DOcZwfLTxtZTb2w
89qeWJa+/m5s43lk/cTfISRULRXZyGi5KsrChPGCZ1n9JjtoXfxF/ZloOhDWCqa6
LjROIOfAhmqoLYPudNdBoNyPafmlinY7SpHtPWbz7ylhZuZbOb7bQNUc016GUiij
aifZUuYU9hB32/4xlhfLqg==
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP15_1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
KYzdjlFdSr2HszvTylDldEFLQ6YBSHkZ1XSRbnrkoecihCdUO1Q7f3kO4OH8ptx9
xQ/eT7vZs3Q34fBI8c6b7akcNy6lzOhemVZ8R4hYloy53kmRDm2DypZ9rjcH9dH/
eZWg3OeCs8ZA+iNictx671oMXwRs0m0v6lQUAhFOkW0mvY6OLe5oOo9/EP2ROWDQ
YB3iQRf+deqcu2X1fILcny5wlNJcgMQTRcKhc2MylBYfXpGfPw0Z5pnup7ItswML
GTJlVw8ReTqo/+1ofDFixA5Gsz9ZjPWlqzWctcKyO4Vy9rKj6sWifrRyESwGmT67
ufQcN5gl+Znq8tquN96yIw==

`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 26560)
`pragma protect data_block
P2Jc/SIiCmWN5vc8h0IS9gS21FwDGzTl3tAqCFS4jSPIAp2xG8cJlbYbLOohkoOB
v3BjyVugC7knTqqjvHgOh1W7/agqUtDwiiuPdbq+ffc3uuD0nJCLhYPdMWQD42+R
ig5ja+2vzVor9N+UldKDDWEo2pjAKUsQWGjta++utjZhPk8H3sHkf/BiJ0pOO0P3
LRormG0L+FOO80zqTactuDLrxtetznAjp30NdE/tBu2n3uTwoBquc2K7GRrQLJzr
99doc1YHUSeaUr7gRoM/N3vXYjvBk+Rzq0yJHpulP1/JuLZXxQL+2LcLN1qmvgVv
vjHmSt4e8/DwrquwUwnsbOOrtB3UAavIJIzgFVeQ3ukv1rttkOQWBBQGRzMyNG2E
MsGTwa2o26iCnZatiJcIqrT4hkAoFpl4glJv07nQY/WaoHHkdP5EUBGi2e5QdUBK
ClCJ7C19OGKs/BBb0zWa3MzswHKjZHrKn9RUQ4t/yihmK/uKCnEsADTcrKEUD3qI
2Zd++SO7YSMaOem3J6tia6nD7vOcOiKRmfSygXWXCtniFlIBWrGk6Y3c4G5Q4hpu
K5E7Jy0GG3cUKPeL+5RiHSQoMOkIHmXTfqo/hHj9UEewA9wum/Zu1ZDPC4T3ePZf
tvNBMiqKA626ZlXrmlxdkKFgXxopFsh1lSfCWToou/GsLkGY85c2wLkCs7a8sGTt
hzo2iJMpy6zMBMf0l9x/SG3Iis7BU+awesalgjkwbJaU47qin3vfW3ee/vVJD4pB
4KXcbzVE+BW1p58+CFNT6AF7PVnuzSIij0eMgjth/df72csIutG4n7C/5RDVYCwl
sVBa6OwPltduRsaGmRlcEU4IYo6ZUURnMnEbzA9Q5TwCTh7S2lIOeUvlQKd6PmGs
tPAn25+QOyH6DqQmK6hWXsywzxFpKGgcstsRHwZGC4p7cANxqSPoDtWE+xYkSf0B
kIOlSDSu4idCtJBGPi+aulhlRDhYM8WlnCLiNq4+WhLtyA9l2PTxSw4L+baMXf7/
u1nC8C70fFeovXKVm7nZfpHLObz9NtT9od/TADgs3Oli+G3nFeH2uYsS/7+G8fG9
tdtgyZbxuVaaXH4rs4vO66UU2gLl31wXTGkcwR4rIjN/7Us6zHT+JsEHNVdb/msS
tDJ1TSlqmMHufMFonHy44veJ1L70kMGNYe2qOOOUsh1EePlixZw5KmN7SR5atTDm
ZH1581IUNpY54bvSMek3y9vwb5dWw3XR3p3TG91ZeUZZtz72PyivP1Q97/1iEoei
akhsHcoFMFXBlSFOTGQyqKaAxoOcsXXJEkhNde636nH0EoqCDRQ8BJxsk9V4DmXc
xVGekf8SAEbX66L4gG7DUpT3BAAF4aoqtFhGHYb3qg3jvoxkhsLVoZvDYrV8oovz
n2ol8Hx7zSGWgrgHzfR5bZRDBU3Fd2UKZyF8/HT2APlrSOKWouTOZ+5MyvETvW7w
pqO8Pxav+tHQhr0taaK//vs1S0B77NBWLCmT9aAkAwM1e+o0ygJN5Xm23ZQNIBuj
ZUvrGrpueRCef9CPrQZDJ0NQFig1VjJTLZvLbNpRaH+mN8VRoWwtmtosxgsoaORQ
4z8bTiHS1QzmKGKnINsLumHQmcaddT2AkDKdT4IQ3ypOYPPPyiEr33Ki8IT5Jnpj
57EwS0O5nigEEsfUk2QxBTwNHfFFuUq/Kn42r4jwCI5BBWLButF7+M7wMeGi5T7I
MqIAr5YdOKY6vMOlLpC3f7nJWkG1d7mTzHTecUYIaCgwqOJTvucwoK+3DHecDfgD
LJPg1rEnug5yEJpu/wFzqYgKAbUGCt/OI2zj3XuOWWTeKw1ncIyvYpFXSwL+oZZ5
KpRjHKL6GG5sRM8UG/wpM5ulpRR9gSmmjRrYu9zOEzBkGJj8bgw6RDERYesRMyeX
ph3L/VGP+GGM+M+uhmOHosb89mqsTeDU89KYXaR8HM6e8ifD0w/wvnLcr8YDFY8q
6XulHde+/igBJY7q8PI2EVgRdPFl1ltLSuOr4u+0WMy8JDKJU8XZJGm9NJI775Qi
pfFecseQSy79efhqlJJstbLQGOA/VQYx/s4QofgZJZncdC4ORiYrthF6DWWfSpHl
5AW0VHl65WcwDd8ByWnAQnk/MzZDSoXL2sDgY4GpfJ7FtqNP921l6CcmDm9e9YHO
bWIZ6amHvSWsqaFrx7b36QUEPWYe/K7Dig5Da000vBV03I3AQExZHFU3cdus2GdL
v8/FQNrQSoseaiyR0VRxsh07cTEpZgHenYOdiW3f+nSP1/brlMG4rzpxDX7Sez62
/PmEJgeUky5hFVqiKHaAXOMjc86G3tyzPy+R9m8xHChe8pnUovboUsYJ9gt4KWO9
g8PXxnbgVW7p4UoGi0rHHRhu15Gd/e+8c4iWlOcG3FizZrccPMY7S+hGx5dz9gQw
RSfyvQe2ajeOCbu6nxsWU8o98D+aQQMl4NFFRUZaVdoF7OdQ1C7e04S5n2amHHof
1fQZ1o/+OTbeTeCZEq8xXT9RmHYbhNcUmWe2ZjyI283yIB/HDTsWHtB4bd+Mt/G7
m6X3nAm4L5Gtph1eBsvki+YGus04mhH0D60IYxBhAPhflfWo5rKpoW7YV012CLcD
ahlxpULPRpVdoJUTiUNIQjtw9OYN30Fv89NPz/5KwfVichjPYOpAP14DbsdLIXT1
M0qi2CZKjbMbRVGLuwfQamKNqdqS+ZYCzO+QHgmwDhGIU3U7BxgZ48W25KD9AR5a
OpNBtI4jOFkYKDfAIzd7hmmhk6hV68OfgQrO/nOLVWds7tVMgCWWCZugGw9s+SFB
F8fbLlnMHa4MPjI/Ew9USLN6CiSdENRsbjSATesNye+IajgVb9IorDWX1Qp+tF4s
GeYc3UXs3DtF9H58wCBy1oU7u9QfMlLaj4udSoQX/RNBBSHMQLzMREYq4K65uoq9
AnVvqRjUQPEdOlRhM8AcGTYG7O57U5uLqMlC8ZYoqEzBweh0bzkL7lgzhW2KZ8ia
BWeZNNILKXUOE8/p0qhtxeqn6mKFuzFBMftVv7/6YmP6u5M5MJsYIGz/ppcG4TLQ
907Wzjb5UNririybgo4gfAHYmxIeK/CBysEJxA52bZTgNsNXzFh48U1hSMGPoesa
PcIvenv68YQEIvq5JQGLdDF1hkD4hspP3MPPh3j8QSDySwbyOWQx5W6JdM7xkAoo
uN4yO+WIS7tOz/3dElKMJx9Fw9AH4t8ZMyW82RTsL0rU6tZczbrhaY704IXI3gLy
8a7Xj3tc+N/2humLcyASsAhVFrC18sLh7nV0Zc/zPABDzxsqD+aJiZH7SBIzcbYn
TmW0Ru8WLtOQmOYlAtrSzMEiHSY1sdvxyjrH0zWNd3ZIOOdG8Hk8IgGsD5tCCXpW
5hvC6AfZola9RA79Ngf1zKEHnlfCxrnvB7DG1+M+sgp1doRt9CiHBlHwV2QomYhA
y5m4cSIGulU2qB9wexskMUKcjkP3nZAeBBiA3pAvNvUUmvy0TI2Azt8d+0fyGmyw
DgP817fR+7SvziYeMANNpP9yxILTgf0/qa5ivmprms92WBR/kO58vmbQ+P6OltA3
h2BehnanoVeWA87lLi4jti2tnx+JT207YVYI8y4XdBdwrv0Zxu8qwPPjNt6Efber
lPyFyOZIZI8lb0u8ZJm6rPixa/f6/HO2LiisDdOAtuMzvYDksKBCjV15cRSCVVj+
KnsbiSkfuvOlEXWAypIf0UszpNLOKotR2lk2kilHUxTpU71X5zOUX7SvYme4ihl1
p5PunydAt5ax+ercedQAq9oZePQ1N7Ngyv1/xwqK1gIxvt+0FMUiGKxwBlhOCN6M
67G4KU7Asl6zsgSgPKEOT7kLGva9nt1098HSuorWHjAcb0rAG4fzIEFbRQo15qAV
5JBj2Bu9Z2rs1HeuiFWymOE3jE+032gCEp5Nozgj8S66mt9P64jKAunvZyT0Qxh+
BRuaMt3z7mXj8vt65GaTdBUMrzDI8qlsNJZ0KulcYYLjc3NBZ6mFaT6GbBgMLCWA
Ao3IEzLWEgg/Uwdtoe5Jxh6QOuEyec8d/nvADqfSErQF93WAjj5Zp9QGX9LzCCKh
VKLWF3GTEvAvu/6/J4MKkRzott/WfJMyFtPJO5ncA6aK5i0+ALnnOD9VrTkAL4/R
SrGgj3c/POltfA9ZiBek5m3loJp6T3T7/MsJno71grhpP5l6o6LcBdiN9D1gVRJn
8NwunA2zauw9wtSUKpjlvY/ngVtaaSLSqfqZfwOZ+GhRrsFReiuEDhFrqco055L7
mlV487PBCsuEBoJ1W4136nxpU/kVhry/ooxzlHKpGdVJcd88OQ8QrOHxH2TahoRQ
/C6Alm+Zdsb7Qr8Hk/LokIFs15EULQ4E4N5mRzIpaPFm9o24evEglnXYRx/i2VOC
U/Ss+3HHjHovGNXHK5oFjFdZj9W9TrDiT0X/3zeLW0Eu2MRK5WqDy0enqQpzUMl8
mpEiEKpn1/kQEahmFEW3e8f8TUjW8rB/nq29QgeU41qGBQTZdcYJ85pPLYPTaUyq
/3RISTprGBagQRvuuWUoVdKUb4e1LcFvPn0BxZAu35oT0VwHTDAqqZ6jhakHPENR
DJelHAfTc59KqKTlGzYT9hQyYhTWIFORQlCVQ8P1E9PC8BAdpY59kzulW4Ekg25B
ZmXBtMsiWQ9sw9zHd03O+CYIitHJ4eTQZRw+DDBJKL5YfG1Z5vCcq5oAaPq3x9iH
uXJlOOfqLJPg967rXyOCmYxMnm1eIyYITRCuKZKylohqQgL5dfMvt+He6eIPQZxG
PWUDPpRRhB6ydTXkwJRXU8okQowYyYLnwouck2qdi6v4JC56Tqa7OjlhWMWvD6dw
7HfSsrYQSR6Ae8/iWUZEm7smIJy1sarwmkkFfzCWC01u+zw2xyCV9VXe7NrbkZWI
wYQslMYns5ZY4mS+3pjWtWQl3A9Kt4x65R91NxRMTrwazkF6ps4GgEy5X6eP53gM
BEFRJmqdK4aHriAbqXvPapuEI+2pt+AYsoEvTTPhP/FLIkOienuJEt7zhB+g+DIT
1RhiGJMsfeNhPOzy4zaTD7+/4CPftQV0jJFZGy5gDVRyDU8wKh7xKw4wWHvzwxvW
rpKNX99EpOhWkU257CIGoTBUGiP+qqDcVmwFYOxJUWxe0r3HEhgCqRBJEHGrptTs
TiqLJwcDLIfgq8bmaH06H6ZNk5XZQmmJPS1gCxfJ3IH5H+7J8lAXj+5SLR6+RuwV
6cvMU+Kh/jVHPGLsXcmfzrnA/OxjpjB149y2k+IzhRydHgWA8Mef+pxmyxlN9oXB
PVECqpVPYX27TqWcpVDPp2bBfJEYrfX9dsO3IXRIhqCcT99U4tvVOhGfaydbQsVq
l3GWlI3HxRqSjCZoSx1eRA5QMjKuBniKThNE0Krm4dn+5GC8SEnfXMG3bDukc2mx
kPRARXiY8WFX9onjAfY8JfDLJQQkpKPc6+BCafQ1zjl9A2j3tW19KNWibh7vpJEa
IYpmsk7BdyeDyiVQXFh/6T4+uhwcHPlAFwh/e63dsqOZHWbameMy1rZJrtRNIkKk
fztWJw0y9+a35jWLbjmcnQVTfYh+OH6C/yx+58BgFM1klxfhZ0vUxWVK3BH7nJe7
tIoSFRDdnam1RgPE7HKZ6JqQoHS+s8z8HupC1CdBzGpPw0Vbh07jNvmBo+l89MMa
eq4NJF7IsRy/M6pNZ0K1X70tiMzXkEFMgElJcgjY9pAQCFe/yxI456ML4ucRcaWx
O2IEjX9CHwqvy0HvWY0qnELTIuS6tylqK1pjQR1ni2t0rb3IyiF11xAY9yc3WZHB
wcrIa1BtfyIVGs9T250Rxw12KikoJzeCjUDVu42NOv8jefrwDwqNRrYTiuJzryyQ
NWJ9G9zxf04daIbyx7z+ITSdmS5jlI3Gvp7EMsxYUX6yzHdiC7Kpt9WaD0mMu3v2
DBG7IiX2YuDBXnA67Cls0jbyBXYJY0mc5KXUdl90melgmwqsIsnMTDuejyDDF+wS
HhRhCtrsJkr5UMtjp0jybcErCCttgOBRjYkvT3feuCVuwqEwUvxJHX0bbFF/M223
QoLqRGItWP+qjC2Cj3Csk7SVHg2ACwyGrW8KL61OeXKyAjbfoAOWuGT6ygczV3B3
oNsVvi2fKSfkpWcpGE18cbEztHSTZCAT0NVQEddXAEIty1evMNm55y9pry8mfY/I
wo4nJoHMcfwYMd5uXe64xFRn2UKev44NfupRiSV9N79u7JlgD4OZlBWHrkALxStK
Uwu8qLsRmVVCIeDUiZb6DbJAospHeMsT2KgjKdZdfsmDmqFSA1+jtir5MbiVJJRP
vxmdif2Fq1Wr7JXTbpuhpAl09dA0VIuYP/Il1I0q2DxUMLyIVZsx5CrpiddiK8gA
DBELOPQA6x6Xs5OJiAR5L7UZA2umFIFkHblH4ioOjC4FEK+ls+09+eOrYXyQzdZ5
Sqb7x/NUyMPKsK3nhlhIC6DIu8kJlAeziYaGv2J4H6hQVteqL6i71DTss8YXsLud
3laP0JPGW6k1ogkxFoWMjFbQAjUJwyBKND+AHfRKIaMiTPlwJZ+oK0Bkl2+aI1Ud
U2LRASNcZN1Qqd5wk06fiehO9hASkicniEeEPZtB9nOxRawk6/g54JAZ0+hyuXRG
iPFmcb9DUxwFybu55l+6z9KZksCq5YRIRA3NEqWj0mCunaLz7paYYXPmmXbvdJ/B
NTX2ycEAqdhvzA7wrCKRTET+CPeCFg0fpKqG28Z1RtQL/+LNO3ScqcbCVfKE5iQZ
SWE0JMTPjuvrPal9syuAXxgwzJl0fwn6Hrc4ekc5aXKDOh431Dg9kdzZc6oEMzVu
PiFt7fFoI+Cg0EhW+oDp64MoEZ/m/0kNdIKV9wD3KaGFHH4NJOGWDWlE30hy4I33
I8vl9xl0cCdubwBH2wBlHXoFun2HFahK+Z29jWNjaA6M8/ottFNYtP0yToCKywTo
0u8qgVTVs3Fy+tRVmRH0EOL5KJrEBQ10t1imgcDcpjsuHC2vU3YzuGj1Zm7ZgctX
RgVr45v7FSR9myRHp7VGujrin9v0TMGgDt2X9KE6vAK9tLcgDXsX59MR8w4X9I51
HwAj9MCNm9f5iWvbsKpeNm10nr62k6DVBUXCtdj35oiKxz3CVz7FlYRK8bK6n1Ck
Y6FSoHItluvdPLDPvm9h8x5a+Q7YSPfOPzmD4HgBxYkgDluBS9Lg7iiVyp/LWqdW
l70YPVwVhPhBWDgMFPmHxj93DkKctZexGZu2A0eEKPO94CyUvogWtoRdWl0LndoU
5FPggJWCDRpAS7PnJ7FLkwdXTqGmDdN2tpP9xo8ikSXTUgoTqgrWX21iwlM9n1P4
AaNtugYMhnlEfh9ECMjjwqrr2V2m8AEfFEUzGTR6fJkNjAFv/HiZmFnL/hOJU5aI
milddqeSo7ATDrY9JR2hVJKyD81wC8Sd29o0Td3UQK9jPqWjXWVmC7b6ZLHs2jfw
BIZVD7imG2tZIAvEflIMVKvdABgPDR9EnqK5gShIfFL8+ab7v/j0zgZ8RYyxwEGK
nft5b0NeqOqK9T/0vk8Xpx2TojfAv4O5X6YbOHzbRIZHiILUVunH12H2VCoMCjwl
2YIQt1qjsvGt1B0K+ZlHTgoc/TBUZkPYtT0oMegLOfrA8Is++hg37pYem9obxaMG
RBylx//wDBZSX6+UTlQWdq7RumY86p4vsmn98LeK6SXCouUHWN37A+7vOG1fEvJ9
KTtZFVLoz0H0iAuYSK3iesi+vI7jklC+i3UIJmJcO2o9cAiDzROjewE+QXzXjL7K
4JtUDM2wKbSoNf/mrEGnWFsfvts3rywB0lcBuQBpPh7uBjoGguHCSM/ijU1dZ5A/
nV5q8EXpnSXMDeB6VIDuqXa0WrgTJChslcCyfRbOenJMxM2nFcJkzGBjjdENlWUc
hipNk0SksD1pW2y1K6yyNZaEDi1dEoL5klrZ3zGQVhSbLalf8lljr+PjSsV+HqI6
Y4xYh6I+atLix/83B30rHlTc8iRhZ1K63IY7zAuMorU/onTj9XGgfEo64fS3vrDA
CPYagREyhDS5vsl3prstHpYSExtcnG0cZUStocxupwLUNjqJSZBSi4nirfQsKZft
WJgjBJAB9HEmtshXzGNcvKzHe82d8X1XP//P8HUDXOdY/DfVmWOv/ZACRGUuXvme
KV+IedHhtUHxTKDLyTOzDRhLrKs2oRFvzSTGYBd4wBgd1i3KEDbs9iv0vPOvPm+f
nDsR15SDuc/vSvElqYPHHJVU7Nt6gNo3Jv3OcSzrOfB06fAiaWI2H0u2pB2q7+Wb
hfZr6i0Y6j6Q3QZZ4/4GPxUsGEzBdv/4R40RlFU7l5Bkwn/mTQB7QwYxRi9l540k
uR2hbL3a0NnELNghgA0wGF65CcOeV4WZjyLe5yaZcH5kLuYMx+3nFIpTQ6GzO8kk
7iOecGiLzzbt4LbPQ0DCzjnf7fAURRjvPZkWEiIRZwBlBP4Z2slxqnJQ7Byhqk3N
nIs3CRhL9eZ12sVeYn+aOizW8B7YCvQg5mYREQ7e/QhttG6ZieAz8GH1zk1wNf8R
L7usR3/0vpmepACu9DOvkf5Etqn7DeqbivgN8l+xyEMrZpAXtWD2rSWOev1s1QgE
28KUY8CNi9TK77elUUuU8rcbQaXzLpdl/GB5ErgkDnOr1zukUwSCHpEWSswNyZ3C
qlFoHFOLX+VP8XhGmzN4OgTEe10CIlkxtCFoQZXi44XrcmoWRwL7qeXyQ/GZhSzO
yFgIEAiozr/MsV6qnBYJYFGW+KtNNoL6qRGd85FnoU1zqYPHV7mDVooOg09a3Cdu
nj3iZfoZx82w2N6ulNai92j2d1Q8hXR3X9Ce05La413wUwJk/9po2sS7Aa931StI
qO+D7+TFBvJD4ATp40eQifZUSM0VSHEeyG4KQGcXew5T7VMMSJ4kDIbd1nT+Z611
/v0j8ab44xKHkCX7UmEO52g8p0PIC8eaEJ4IX+q6doJx0VI/jkKdCqjSXQVwAtK4
xz/zwb5U0gQcX6AIXnwxykfIWS7quCdCKux1PBFrsuz2XPjzBon7mrmPnYH42aLF
Mm7OhzJ34fMcclmEACPM9SHJNTublCgkSXYK41w9rX/x9ltV5y2OFDNccQEcHWFX
snHjW8Y7kucaXn/ewyjabrvUTzTk8tL0RQprNicZtoD0bvL++WrvSCJF3HzvWwZY
MKn4PjpvgzT6CzdiQ9ySzrCIxznqoXB8pWBpywYHIfAt2SNCi7sx00ayCRhhPZXi
2OGVp3CvXtxrEfOfNWseMzJl7087cwpUcVdDF+pRQuZWiZQe0/3OyOZAku13rsQ6
KJvpKyE0cBkT2OkT8VfLX3jSTjVhCkJdGTLl9TAIQbBADM/ApnSe10eK8MnS8dG3
X37inX9vaTpwE/if/wKEn0MhDXAlf/7nSZVwggr5vR6i4hpqrlxDqw9z3tiDTfIX
PdLr/7cDp/ABKQ9OddOQr/mmtGya/lo3HQ/Pbj5x+tGdL5BuZdHlJPtldvoT7ujr
KQxU2EsOo7ar5VcnCvuH9CM41rp0AMDCIirxvqLfyodCK/9QNWRtiMFShzSxG2e4
OX0eLyOyWig3ssni25T3ApCG/0fMhalS7NPHN9vIxLZB44808twSNT88SQLASD+R
frlWx9t9gCarqAvkgnVLtTFoypCP0HWTHPqnk190wXY17DmTpDutLaLU/cpCd3pf
LU3aNHWr8EWsuNSf+1TzVGJhJyaMVR5OrM0pXScqNoBCooR27kZXKdCsqaLephhL
srX9czipCYOxDmqqx0XeaVMkOyiHnfdJiiWkd9lXjdo7cNvHG1e0BUv3tnt7BK/q
tOhmMqM3ldD+2pJmvAocWRMfDEdPKazUJ7l4veGqkn59YDSbvsdIL0mYZ6pN5/85
qzuAfG+Y3D2uelyEhzMs56rvt/509lRAX2QRID7EyKfkRP78WpaWCNsLmrpeCskM
pkZFwiS6bcl2RxlL16A3O73JGpq4Lh3QZnq3+tzwv8YrVu30yIhk3AHVY323gzFq
Tvc7lEkmha8TWZEg7zOBeoy7E3OTjNYHdv16hTfCaarVUTCT7biTmrT71yhZLsRV
kkWNtWP7ogqPlX7CcqkrRTZoWyvsSkmwN5ApHUfEqhC9eQwVZGyeSGTXFRz1q+GK
DEhWiT544f30XI2JTouNCfCtiTnYxSqTSi7PP0EYB34mHl3wfzvCCHNcUvietWMX
CQivf+VPS7r8ErAUwVsQ/lnJF0W2TcbcFgXjsEVi0jbfziGyDs8xXNlpPBrXEF01
ycR/6c+nDSSz/11yQzCgSxW6gbtpRbAllyIlE71SjkitYI8D716HhmxFq3GvoHii
bnGrGyE3jruUFA/tpiwvX4Lgw6N43oOXkg4lGGX4AC8E+5Chr/jArC9vr9Z7by5I
DqKUL8Z4yPHUL3K89PsAFqWPNUk3QIGGCeXIOVNqAys4Hi2RdRLZ1b+p7kmcn55S
77jVk2X4FA4pHUMRMIcH0KppMp/qztqnWy4GUYz/xBhW/9+iAPDrd7YBM3dg8VEP
YYVS+GX3Aehg7feLShNQ3Qio6R+qhk27OhOdKIjgvbjG3n+dw7a9PMCvzvmhUcdp
ARx1RBoXI7xL6H2gihCDWi520EBZLyVgMRC2Ea6fVTNPwwLvr2PVzkYNuRxdLvz3
2pDe0s4Nd/767p9EgSqvbfkfZsEVr7L56yWrkr9+55kRKqfFEvSgP9e3+tduR0qT
aiK+4sITRlkctCOOv06nZPbu708CMvS4tFjUJrzUMEGL4/BKjFSOmIWrEQXqm70U
GEFE4RYlV8hMaaLoZst/A6IidZqr+3Bdf/BgHzummtTnqJLx5oOcGIOTrvFe73os
PRwIeDDQLZBCI4ErdM019haW6UGz49cXY4zsDjglmnQiVthrWT082+Dt/eeswaly
IbU1p/bmfuFe7INn3SmRqqVpIbGsdSWbUZAodOJV2na7KCIWOaQ/XIEP+wpK7Yda
ZK6g9zQiEhkw027FejBtJdfkCvS1LEgfzlrhcZbSvSisqIuBn6faXv835ZvRLWdF
ezXpZYs9jsaTAx93x1XEzG6S7vdM4/panHKpHb11ptHoscKbhXcrhdB+0hL8VcgO
7rVRPam4giW1GAsT0f6e8wC7bY7yzI/7yjIjaZc4mFj8u4VCKe/z81s09yqXgU9K
0C8GkOFLYoAMy4SrSR2aUFiN17lgUkEI5nwM5eYlF3EHlJKK2B/LDAyLyO2GQaCn
l6hJTwxsNfTChzjG0LNGw/xUoM9guBZ2YeiETcSlIhZsRC5WzC4ELRlLMaPf2dyg
IcZ+u2pz8IrsszFCVrXrX+WOZ2OsOi7dnGLED6HTsYbZ1nOamqEM7d/2arzkGKgv
/4VVa194YLuUC8gxtd50mW6NWtBaVFwT+J6tgpQe9kIVGjabCtSgLKd6Igh7weaf
vfWh1gVyYWAJTuCpg/aE6Qx1ipN9yRgqran0hEHcx+G1oMG1td4E0MTamgvXT+C3
XJ/0EEclCs9aueYNP1TX3qtkySBMIG7GOWbDC2CvHuLIW2szaX5laPTtY1CZNUTa
X1pnE1muFnu+UDrq+a2EOsZGGGh0rtvQ3QXxf1NinAGAV0VYQoy6adyCPQUnf/mz
NsLRjtgEnCeD6zbNRB/r3HBDogOeiT/6SO9a6yAdV2h4PaKXYfx58hvNR+gxgsyO
Ln2GMANnofZdxHi1YLCQd6M3Vmqf33g1S0VdUzIyAyt4iAc5zk2kyB0lMVMFFu5S
v5JUP0veLZHFRrzxYocwPRtEVUjLfzUnOY3SgRvs9Vdm3Hm8wJ9vjvF3T40rjusT
oGMW7UC9j2kC1KVK/IIaiIahQI5yZjEz14IqsFLKeEuNF8m88ztNGPSG0qFkvfB7
/G5rDB4QY74bEpUvg6ZrQs+ykuRCA/VovpntZiYPJlHpYhPLjYP5sbHP6+WZoHiF
+AJS1r/Djg7aFQjglXdAxgOt8l0XSU5FWlkXB8QYKj6w+GXCo8vF0A72S9Ilab/u
L1OZOwgV4Qb3biGsnORksl2mI8t5jBLcV01spb2DROeoKjW0F2t2wI8arQy7WRRH
9BEg1iKRyenRDtjEwyIv+83LnfN/0l7c3uKhDD86a42IPfE4b+S8IvTWFkryMmoM
kxH81pdipLuEzlA/GgUvtQRx3XVlHVp/lL/0YFyvafDBT1K0RJ/ioV2MymVG9fKw
Mlf8lHw1LcW9o+4Umbo/F2P/hUBfbOoWQFCkwt/xkbYVScHQw9/vUqTr3OYGAKo4
Xyt7oI70xNLkmESJSY0WvrqVGCiinN73CydCJ6FzJcvVQgpvyxAc/c9ok3A0hDNo
q3ecDVHkMEUH1Dc9bIaWXU7wkWj75FO+bjGmAyuuPJekWuCAls1MwNj9xg4i9T1Q
jKFVvKbf3E60HWyyoWbsTyseFvtNSlpGk+TbQzSGOt23Bj+fn2dN2tDeeh+c+lH3
dhgfGe0xW5fkwDQdUah0LSgPRyXD/beCK9TXPeQ0fzyBPv5vohhTz5mBNqvYBwD5
RArl4xf2FEY2PZvFQCr7/F/7izDnuIOpQ6Myaz4HUtjDzAaMmvEWqIlr28DUHXJi
UlR/B5bj6KIUOt+OWDSPtMYuLG0Gt6/Q0lQSAy8CLV51g7ty2CoEo2N/rBZlT75x
X82SHIJ2j8Sz0XiU5X08YFX9RaMthG/A0/D8t+saJ5RX18SX/qIhhOdxs33X2SRW
kqyNo5XtK1ISBv34s+t3NxwTTns8XCzFPDMvYvogNWEuEjOHEDd4jOCQPE63Trpp
nt41eke5FavqWE7arYcIM4n8oTUkMvmMUQX9nAR4Y9gV7ZlOS+sSrVIRJwcgbYzM
v75jwHMpdF5v/9H3b8YYUolZNS5CyVV0OVeGB9SeO3WVEDoKQCQvvTNnfJ9DkkDh
nVKH9b/9TUaUzNSjoGMClw462rcTVX6lpLLBdgWU2Wpv8MMry35IkFFgtHGJyXxo
KKdl1iaVdVUS/rYXCul+jX4hwNzr/QtkfqP6mrG8S15mOzJeT9gyd4h3SgKNVrRV
yuj/lvcmI5oSIlqLAbtyJp54UIk2oAV6E3aiIFQv+6nXC4AUhFbqkLrZ/zNEksUP
lpM/HzURSYbFbGwGCGJA/DJ2K+qkPT6V7F/IxCW0sAcbx/MVrYUdRed3ofQ6ldoM
G4Jj2A7xfjJsSHtsiWS8Qf4mIrwqDTiAJ59MP7FTXgw4QwBsYhyJlBt7AQyfp8b9
dO+2H2O4xGvDTyrTuynlVCV9CRFWooX6KeJuKbPBVO1ms2z7DGXbWpLbc+imeCJg
S9Aj8RtNp3R/X4ewnURi57cdOe7kXaqEirL0x5bmzOoUig5bFRrbx1m18KErkToX
G1t1y2/lvmf6CT0CcpuOU2amd9gs4I8+YM0gs9hsCLP9JNd5cPmlWmeaGzaObNBD
iMneaFiWycaVee27Q3Wls9AZEOQhzk551Rw87c7C/jrKOWRpjSAvhupR6pGdpfdp
enK9gdCKZSK3+b32mOb09Zp7a5op6JqI7kNM/vRYXsoLb014p81qN0BZ/gyzvghD
FWU44rgrhICOwrwI34daYZQ0AST5AUc3g4m+7w42AH6CccFN/sY5HFGclenBuUnC
kPhOFRMmy5F6xk0C6UV3RDMhAZFG0nJRm5nB14w7NXm+CPQutooJZ06wpfGKGDJ0
vEdHOLpRECK05rQfc2lfG1JMtVGLlOo8IbhQh9lgCvfj5AdB1iw7I9KLIhmKq9n9
x9jbFcUtOLxN4pkuy3S2Y3MPB/epjWX9nETT+LE/PithQRcU1FYpN1RKCQ7P6elG
SAAxMa6G1DJiEjn7FG26YOdBNuwcyCmgW6u/RpEkCRyDtgKlxad4s5DDOIrHyE2M
kJzqu0TUPwTALQYBqCMgvCwF7NpKG7xHDfpeXcnk4NtEJxgg/uFX6vtO7ht3r9Rq
hvrZioU0u/K1vbN5gEIt9mVQiljg0WZ8n88DgBONzqKgVRJ6iSiSxZgpCib8uYrE
QN3PavOZmPAfKO61TpfgJYhMCy9h0s+44GV44+3Vn9AGSz2GeOYsdaqrMNhi4zb7
E03eCcqsFQxSwpCTEv/JA/vBxtkoii27GcxwPqHjcpyJ1B3GuWEwBPHNeJXeGZa9
oImShySZu5hLXEJtPYOg4JiaMBSUyJtk2LSY8528FyrgglvCz/UiNtcDdFjg9tNT
nma0VKMIkppclEyL0h1zKedTCmnkJHFMp0xM9Leyo6VWC5C1DSpMPcV5kNGs2yOY
GTo+ROmdHTQF6K+jEm4rYsN9pnzRwJY5HntBsgfnaaCFIBaTPXQEj6R2utXwKAKs
yXhJHw/nActfAjKOAAo4FIlmJz3sLC9IKkKTxO4ckgENcB3ygQ+whK5baA14hnbq
dGoJvkRI48mNwZdsyYNn2GJZ3qdSI/CNJYMAFGgZZZib212WwpwNG6cRb434/My2
BE+zm89aQqnRr7ANdcvdQl02y/s8b4IUvpzTeJwn4MeVNm9GlHDCjH3n5AqI0jsC
aPQ51OA4MoBcswzXK0qLWefAZfvPR/cbv3yANLkRWfTMxO4p3hT84bTIjfCbMtvP
Fcu2OKI8yPCQ/b7Nmr5jxIILwO7RSwqNwmiGBft+6+J8MwWDQJ2899vFr/+7GU/R
TNZBN3dztdel4/SVXodvrRGdfjaETZbUtz30jfGYfzQvXNJS6b+K57Q1XmNzZgeI
IO+k4z1WZ8oZwWhj9ZikRwcJDphUYc+hDhJ0esql1yuM5mwbwj2fddouyW8UfU+n
1b8Z89bpLth3Oje6cQg55/yQxcir4tUa5qQNC2NLQb2mXgwiOJw5TkrgAZgL6lMK
bCC2Sk/t6ySrkMH0/0sFxkCSTCl4ll0nldSY7rPojxCSm6axj0AgI2UaLhHDP2rj
g+/+dhcgfIz3a9wTl3MHm8DyUKHdI7I1gJco3bILrgFqvjvf8RNsUzBdzeomzUsH
hweUHPKA7Yub/glx2SsV7OprnejZ8G7iurs8phjqEP96tAwh20ZH8qSeT9ssiMGx
yqvAjoRJH2pyc/YxMty/rueWpSWzfi/rnQnV6MpKXX0Pdyphs+A67cVXh3cE8j/x
JoypRm27NOzQZfTCYeKQbPW40SApMXVIF74UghNGgcldboLCzZMbHVyvrqF46Ck2
AQIy1zjfYDdeXk85IZRFzuPg6LykI3fC6t12mfnWBJSpg3dFBMfC0y+IX0BDAFgO
+LIAYvlNxpDHNp2nN5npNWB5BYZoPQ6bnwQAxrLb5iVjoas/7jGrPlQtcmhvICuk
iWu3J1Qby2S9rdOzQLUwK3zfYCL7xnO1Ody7WovbwCeKxjXwoaYZrXizzKDiD/Ij
PAhEJBwHtFkeGtDkKAfFuq5J792ZEi7+cWxk8sEdllvjv2LAnBfJB2VRCyH64G6M
OKe2Eba7wDPuUqhZaiZ3hQ+EHoGv6J2nv/4fBByE5x/jRFCvGMBi+sxj0RGTYIR2
l38upnZv7HLgqbC9td218urfpFXYpBmANzgXDlzC7krG8pCopC3Yu1fj0lBgWhIM
ODBfqyXZQ0dPfWDzdR46u/1TWriF0DA3R+bv5iUUAGkJfxAliTOnaVBKJF+vPfqs
Qm/VbzkY+e63gHujF3x5E75fas6EWZVOc/GE2FjlkmjA9oM6HabNaIuVvujmz1Za
l+bpyXUvvO8y+xz17jrQze79/9H7YLJHLHGkn6Ne5wdy+90zvzqjTHVWpI5VdbKQ
gfqYy7zjbG9US5aUUNksUUQUSf8AJcwudj0PvE+EshgryD7KyKH3j3MqaT9y5poY
81KMpa016vCBejioBD/pnMZkMky6DkGcrZEEYcojc7Uvimvhu3RJdtGm3xfcgGmG
a0xG6WW+BtGz83rAuWS9BhRi5jYKPeDXytvbScBOkgM4X+opKhptpvu1Ygwo2O1r
Nc7tSh/1gzvZuPlRBsSuEnx9/zJ6/WSNnyDc13oRyfFgtzJtvJVxBZK9KOa7OJbN
/uQC4Zp25XCTHGUpef+W8xQlCXJ7pty9B+lPITGzvDSqenKtBn46iJ5DLenJGD5s
x1aykqtPCABzKe5IIpvcn08B1MSo3Z2dwYx/GPTxSPIUDeV2BSkyuwcuqi0hhn5B
gRBbh04ZdUd/VFYrYB1qFkzWyv2ZfayY18jL3o7oWK27EMY3rj6y3y0OZKczRa7t
HdltP25u/B8IATM9YEqU5e8QT6zhEBDrIuvPbGit3jcuSVHwZNHg2jvT7aJsA2h7
H+2lrNDHh6pPcEBdecFPufBdYFnSnJ5Zwvasb4YABuEqr5pB/iEpfmKD2JRMO7pc
PucgWZoJMxzosSWABvkXV0il559KWMk2rTA7gsnPnW/m9GappttYij/QMksfVQlG
21bbMqoCjQnVMNCp3tzgAr5GllXckyddV59jld846HhO/1UdaLzB2FagoQU7UGiy
KiklLwqMSo8neiB5q4iCWPlCKTIAdv8H13M/rADhWsaVzlftUjyDY+88IKulgOoO
xKF3Wsth3n1c8Gan04HWlr7sKgj0WPniLLE2rv8pzx6pARcWxBtfTJPgW6c7IBAl
1vSIAJyQhVGVbijmndBz7PBhzpkdKmRGS7ii/imgWrCuTGDMM5IITlK+1CgFBaX0
JoCdg+JtwfLkn+4MmnnpHNwGO67VVNBXIJeLS6Vljvr+pQGLJhRuuj62OGXe0G3C
4HRoNs1WiMbPztsGc3eSwlOHNkrPG64HNgeX1zUcTcNTiGzanSiBVAqxpKODykv4
RmQs0pdxghqs9M9Ugjub/VxY6NeBydURlfWbJBFQNJ5TyXapgHFrqngsP2Hc4vnQ
Tw2NvVbVDEqwVJeZ62RgaG5WOCHdP7hCemiobAH+dXuJ6kIDgtx1k8l+pjUn353t
KWt5UdKc/Yko5Gr0ujue6uuGZJf3f+8TRKz4bvdYhspa8SC+0RtUAoy69Yn+e1XQ
Ar2/OE9t3AouJsuzFmeGyPj7Lp3SNZwO+dNaLt6tYdLZOd/HSYPZi95e1VgwLfjp
p8Dahx44EYA0Br+iuKemyt1OewAgPAKmUxCq4w9Sgau31+4jOrH00aZJ4Hp/CFeq
f9IH1rZA0ZTnQx0FYIAvJgknr8qJSBvkkmeAZl1paqlBQpO+4Ou+FAOhS85aHByX
OdwI58roIiX3FIidCvo8TVZ+513Xm5yiao4uKbHntUZCJtsqn2MWR+o2n/cIPwTD
ApgUh1AxrXp2vr+3N65nEl4UOoTr5gvPN+7niFjLwHMG8IXBL4kzhUrPgBLnpkgs
2sw0BGZgC/sfEtMiTE31PxtgshnTJIpr0v0G2hB081aOchLRtlDDh5NOfx7zmEV1
CrHeV1cfIFtUkDCPhu6ImDhs7sgVexjlNmheNXM5vv2Zly5mHEpkCzUHl+DmFuLs
ZYuWRURH2CeIJJa2knE3n5CX+oTdILSGVUZzkL96tw4vNa1/P8HfBcbIbMzQ5p6b
UK5sRJem5dc4myx1prCfpc8jEN70wwKrV/3EA0oSeRiKMCpvtzIr8Sm7/e2OBSE2
9x9Zekr0xtRNMpHyMWA5DxXQwKZ9HvxbAqPU2jpOajKN1wbiY3/hJJDPiIyQwOY1
sCkXwqhduuWuqZMdybj+rYsQ1DMoSiOpTfpT/5eMw4yMPEJZiCa/lRN1uJdYKZ8O
hkc6GiMpMKCPuuRwSeq5ImwA0cAPCr9zlybGaGzauMdio+l5e8Rm2MBh1J8j24pW
9teesDFoYE/fjG7l7/qWrgAyfwq2StSCuIxvhnKmE8EnL7mik3izKbBDZqW6AEIM
B653kqXFEUlfFcPzDRAhtnggDJw377Uf+glx5c0ZParfA+FNgl34GIXx8bHrUtzH
nCy8CBMNKsk8mXUoNKQAVi3BLBj6tCZP+C/hU4lhd/wT55pWFIDs2CCu3WU5HZmo
e1vE+55m/G2Aow5E8Ouzh23BSpCWbTH94Lm4Nrm2CFHSoCQDgAmk0bGKiUp3Ctzg
du1aq/L18EvvjqQjYSlNb9RSxUFwWQk3gys63EFanDhL+iSp3Syxo4PDOuGdTdR2
juXNbR8T/4fRnGqqmanUga+aJhS1hOzfla1hnZVnbYB/aU8svDYH45BGh0UKPahM
Y+HocHNRxlcdTOxjj4bdeTF4TqcnxdtceCbFvNaqt5Zg33sVDJIK4n19MGdumqvE
KPfmX8ycNY5YI6JMSjbuY4wfNNhkoVQay7NqOXwkayb2m/xyj7dSF78uFg12HYd1
Bw7tOPsNLZp/u9iAQPCHItiTNxC7veoA78lM/diYk6t3xo0Pd8dsm+RZ5FrFEv1v
DSZsx8AEKR5tnpbHWu3NiLirpBJLbk6mUJQJycaxUg+0Yr6sDEBnr1pak0fCRPjJ
n65pwti0kF4oFmLRVs5rpGyvM0Tgnzte6+kF0Rq/p7h1ac6foiNK03K1zwH4/mQN
YOHuxF8G4au2xi5kAKR3ph47p5xC7BWSmBAuTi+wF6XcmlfqZNp0R4A+MFlAooIk
jJjx53h98zsWBwbbKQk6WJgwBuynmbqcG/74qyMNqaj3CdbkonthSZVZqqruoqka
qz6K3ww8UOKBklfeVIsHGmIJuYBNUyi56aSart+sBjLH5SdmTSFC5WLhFbbIQH+R
uZ+gRWCE4IJnLnHaOORhoe0TiA7Zs6BY90CHoqbN5Fuda+El8lD8FsHykBmz7yHr
bEQgx80P3DYLZJB00Quv1iJmC/CVMBrIQwR2urY0CCmeZY1a34gLv0D69sDs9YbJ
u2uii/S/FFJ4uYfdvKtAcM5RkvBwbq6JLteTO9Nr5u/NVOXJMHPiDNQ9yGcZm//G
wrQCXCfL/shcTQ/tmdDI+7cv/oJOkNDRUBWobMrLvOrnT0iTd7qvEqERISyrzCNk
2IgIrsc0YaIdM/C1Q82EgqxsshGXNzh04Wi1+PzMU54UAhJfPluDM3XRbpiN7+kD
SNHexuT/61GmNun6smH8SHsGBb30BJ5dzvk0Pf2XxWBC0IWAILDREXwkcPOyU2FD
JK/sTARKgqhFrX0aIqmoEbhgiGPVDfzCGikCjHoMy2OYFWNYV8ILHhpOw7aZlkm5
ilgjgy1q+FPAweT0koobPpwecEpGWU7aLdAqvrddwUOhQTb0kuka4gBtyjthna27
4M+USSfuXT3Z5i0w1OL/iw1Y/CzzPXX/2OknOVDlB13KWyQTQTcGBkutYOM5szgC
+gBW71Z4H9ikZzeVIzlR6idF6uG9MEnUow8t3EA+i0ITJKNZjnQUgX/FEM311muJ
2zS6a0FaEjA7tBhHqhQNL+lVhOf7dRpGmmWz7w3I4YPDwe10JIpI9Mny94GlHnDT
Rw1ChEavP0wHo9x6IOIU4R5K4KaAHycYv+k6fHzGzlXHHr5LFaA6dzL0jtbyUmhw
Py4loJFb8HvelNYZdrWtaCqodpwcuH5EZX5iPgrZGXf+2jw5nk//KLtXgapo8xWW
CtXjqRHl8Xp7AAYoqhHefL522vg2QSbZroCt3thiBZ2WUUdVLkR39w1+FlZmwGN6
65ETGEu4hrkYrwgEER0N7CXEIrLmjLh8n/NMSuP4DrH6fVC0qKDltqYe82ehmLfy
JgBbDqke7N1pAcT18oZH/rPwUcR7e/jOgC0dxeUNL/2xFdd8QYQ/nz1kSaWwSPwx
GrADX2au+ijJbFwVZrvF2Ofwn8FuziS75G5Tte+JUfp+2FzTW/+jMucmF7pJSv7H
DAychUNjX/Z7VDb+KZelvKMov2n4TxPkr+4Ti98maRIFO9BIfQw4LTeVqxgW50YH
2vAKtq6rACkCJ3TtSjIDCwE8L4k45tAePOcQgAWqDnDgESJsEtrGlq8S+vlolyQL
6yvu50p2J4aiI41fDwD95xn4iRyjEzxC8cNdfQ4CAYVpFMfzI0529Yb6vNQCcztu
r5Q91XOAx8jHfxX+N7gEur95qiA0yRaWbIqbT6bHt8pbABD1+qbMmRZikBwpNPJY
i/nZOtza2TtCTqy8YxrzBju8ijTkouHMvmphDfXu8Z4wkh4jtnDieNV1uWP85szW
+5BzdsgwplDRn9kEsRiSPzyb53oOMJ9UGxGBkcHUF7Nv4EnvoJ/A+pA4B02t5MUI
I3xElZFqsPp0dA/W9FGWPn62obo2evw27aPbN2SfoEaAZI9A5DGM4GuMVHxr/oOV
xd0aVmvhV0zvtnu72Ynx6lYZovzVbRZC7m+tul0eRp53jJvYXwLldQPg7GqX/Q+H
2M5l3mRaWEEMhaX2V+cCDAaQwAjXl3aQONpmAeUkEu/x+S3+911Lb3tBdZe+kber
Db/SOhYLw+ASjRWw9Wad1rooaN1YzGvZoMytLp45UsZ+GJpJe8Ie9v2EFUCHJiQ2
Rb3YBG2lAUbghsux6DCUtOYM/3cEVGXDnrAXkEUZUOUHhHhuYdL1AOWLDL4E8ulR
bZAOqn3cJx4UJI//ZJ6SBp5RnKeQEvBrJQMQ8P99CYf92dVCus7tttQyBV3lbS1Q
CZdL6BtkmL6WIJkbX2T098+XyQlHcCGDYrtdwNxZJVnvHqx8pMw4eX4iniXKO9aX
texG5MZiC+L/xqDOuJeoS14X6ipa+CueZkruUhwHzTLb5DXdl40JikcaPalJn1eD
tLrTMoQyV4TE+VSUqhYFymq8KZN9rGL1RXx8OfY71eJQPjnjD6TmQWskTklE08d2
XCAVUabU7XUxccGjTUuXubAlAfQeX+68gT23tGqyJhFcnpcr18H4c3coiSuBEtX3
Oi1+fnAlLwbK6QaqeJq/9xsu8683/t7GsA6cqiYoIsRJQT1B7MXWtfcH+dQWBERC
C3kfnrn5SwEC3QUKiVkoEbi1ZfmrI5fd3E41YLsKPENjOVjqqV5hdZMaZv8yqIiT
R3DyglsAraA8ZGIQjnChBPBQPIOMHZSJdBzxQpVeEJX97Igzc6QaN6ZENvu76nPU
QItqXDr+LznGKw8AGPkrrOspSP29CPf6LQfpK63SXio23j/Mu6tvznbm7aKgsZIb
unTn3Gkl34L07se6clXVUNTX0k2I85PM1bS55VJYupZaF3//4DPQs/k2eIeKl9o6
KGWQbbaIaM9xbVIv/csLMdNLWK6Xs3KopjEaq6mFcAFvvhsJ+kFladjjwz6Zw9Wd
Ywyi+y5FAFxPRGA/3Cw/dxJjOEimiWzbyggUWwyD/HO0R/PPQ1eSpGT7nUpud2OQ
QpWexo1h9cuSg4y53e8ET+pRgYDZIQWOt8RN+Gzu1uvSfjKVqP251Ar0z5X5hD5k
9z/MNiE4KfWFT521bx5rgxn7UXI2/RS4O60JMl4ShgsW2tm4q5sqhKHeQ+KleltK
sFVtRYosENZ8TcXMtE2huyZeRCHtK5KuGGRtqOhK/IGs/qFs+vPePYndFy9Ox7O2
L1HBD9JgoUvY223VQvW1TTrQKdFf5BJaEdvtaWnHFL5onJY2EZQuuOfUINCWoK8U
ZWn9n4Ba6oHKEPRZRvv+niKRI6SRqc1e1JS7xqMuoPJajvgKQI/9BjeSiI3Clg/z
/FSvpXs/EMwNi6wKQoHlh2CmSgYvjXnyim9feM7e9hKuhMm84cLcJXgTCxAMF5RU
q711Bau7MzVbBsbl4TGamEoYVPK+FlIN+DUtg8weUOdsOON1qfS8WTo6JwURPKLW
x5QjtoZSqTVats3sSOmZPP7po1IN/pyyDrcFTSBZoj7butvymvNL3uyq0NK2ePDp
/0PGoUjACbRPtM3lXSniL8JTFS7POSwz+9fhgsIE0DluYLlUDiRne4dzIALVpRQY
0zpvh01zivYHXGGRd4Z1eElPA+7TmcnCGQ2s3LfJ0898hIULnAKApNbbz02TeEUT
4b9S70SS37T0nPACDjRMTiRzDJojdaTHGc419VjO3La5kKPx/KeVh2Rp5hRzKs/O
MquGgrF1uz+mzAyR7yPMbW7nYw3kcLFeWrPHZILGzdBx4qD2IEOjHHYR8XqA4uH7
Bx0UPwjIAj+UDOkzSAdICXhtH+otAHZJ0sMLQgG0G0pm9leiSbRc1m84y/echI0I
Z9uK6dwpgB8yZ9ufGK/XERS+Of22F+vAPJjDPkfA2oczs/1dfopLE8xA+uTelz3N
ktgmhd2UMajtK439d31BBR8FmsSP0rtKFDFnJoUDgoyvyW1Mt38TcWpdwHwu1dux
LGrQqxYG7ObhGvsKzwWvssNnFZahk7PcrI76T3R9derQMq5O0o7o9y6g+0Vhr1FY
b7MHhJstv/LlIxSE2iwRn7mTaJPJb2FeBpME9+YLwamf/j/wM9+CPD2xPgXq50ji
ZmlYgs90CKsnyZtX2EAm8UESPkwM0/rjhrrDNMSiifq+UFimE6RERiS9z+Faixy1
UZYk7guIxwyf4fGzrHKZGCFCxzvY80ebuEsVdxDqmBFUvxwF2HlGyyD8SyoMTJf4
2To91CyaK//S4L8PLDiBHK2fUmTYnK2C2Y5antPwc2lQjnZjOyB/Nf8WCf2WsPA6
kINMkLiq3CvcOzvVgR5qHbHSQQRatfjTHwMtB1wm/H+5yYf+I/m6fL01H0+J2HX1
CcPuSIIohJOBfBb69aTBwb/j9H+lcDJ2qfMbVRIRHVm3GK3GiglSQjH1uhqCdEQ/
224LGXdR739c4iU307yCxghh6wAwnBaKA7LbE1jwoRlpfuP8xMbDzMisziKQ+3Tg
La48OwEJ9j/eSoUBMBRAjdjMiSFHG5cY0+sfgq44JK+1lEKOcTS/fD89GSIKp0jq
+5GvLEKHlI8ym8PbUUq74vlW9FQP+IGjU3eAKwjxRrqwLiEZF7usm/KxZJJeUNWt
T4nmGCFKBVn+A9dPFaMI49wnI/fhChzrJdowmgLrKRnzXTHYN6+bRv9mOuo+H0zj
pp+EH2WT31fREqH/zJt767xlCA2pBJ0WjnRbAjmgvZHgh1V2/DWaC9XcsvRCDZXa
a5ITt9aqHaCNM+gbr5PgrTaP9bGgbVoq085q1WVoHGdZYfs1ODEu8jgIvjQK9/Nt
89NtZXHcznu6TPn3QSUkaeui1ok27EYmvON0Nn+4WeLC70NCFOTmaB566+fVjxjn
TL9sd85n0+PluuDR7zOESWgG8+VnEnKlZu2PjhPsL5rMCBOTbpKKBmGHoi2SX6Jz
GUq94tE//fnKPPyUnDJKWDU3ojrcwPirvNgceSFwz04zl622+JdZpo988rG9pCjT
BlAALSmPdDwh1Xy4cYWLNDZYOb4Hga8Gty7s0Rf03jp6UEpF2zStH594h0Revy0h
ZEvlAYmkZMBgo6J/xW1J5R6BBDynMT0yQo4z+LoocnmcXfpe63enUIQLLfcFBT61
AL59OV9mubSDVFuhJnX90N7TQYocSRVlBMTJe5nmEeivcD7IyUKU3hPqYB/jtgU7
XdZ2JqXMtQIx3XPxN1E2KbKYS+gi6q2gXb12RjrekpUIIq3Cx3hElqfC7AsvWyHT
cNa2SlgP7B6GbMhqDxQA31m3clo85o0njVIQwj4ezrKQSOsaqMqgHItDmGPoXzy2
sx0WD+lYS/unjHowhMzoZ6aVb78Bwxw6qxpNGqOF+J8NDN0Vg8W8eDeVOzEVvebA
urUtCM2eRBVYECvHIOCAOgpj9T49+9SAabv+jKqCUrqLfVXZH8mcF23ccIeCUcSx
3AE0d+E/8db9pcbuTK5XuBU7EiliN0UCVT1CCd3TcJ1P4aI/RWzhJyXLtE+GBlba
mok/nS5FiP3zQsT/sIC7DYxCEw57D4AmUjL+80XfiHNY8q0agLT+lt8J51UbCRKm
lmaTUDyNHtOtotk1Bn2VeCF/+7/ZtIeG0eEqDb9d0pNlrsw/+zMrRAf+ly/5xblh
pJEQsnT06f14JFbpK1qtzTg4QOY4ukrD5L2VIgzjybcztDdY+Lh1a9yDdpJp7Omt
ShP1MT1yXqa6WEGa5e65IhQrEKOytlLmIqWYq3f7mZB8BM0A2rT5s5qtMORM2kDE
RFNPfsvYA/aPom5gvhutyvAgdkSfGgze3Q8E2hTWnRsgZT1Y+g161PCLVV6DBmnP
lV1NMowW4YUC0qBqeZhwaLzEboEcC1xPcRq5Jz8RI7v02HX4rtMM7RYBAsuVJpjW
CYMoVbeUOhPKEDIwaeGvuminhZ52tA7oSSvTB86ndCiotE3c4dZ6Vjt5K+OYdh1n
xYsIpJzZT5VvKTTl2QDjJj5nI2AQlEOuGeXvjrizsOOWvYPmrd+CgM4arimKkl9I
LTxHHeWrz0j8BOcj6YFqpNRcRTzw7ieUHGTtVlAcsqTHiw4zp9L4O7nepZGvHe04
1vNufgUWbcokaQMddeyXEsV5MvUkIkCdG93q1P5MwiFSD+CEtYID6s1Hm4uG584k
Em51joD4MkEBemONDJsLrpQ2U+I9ppGWtQxu6Yu0bu/1pM4h8+0chm55PHvxLD9Y
ZiAcxqPfo+Kqwz5AliiB/tING3ULcoLdUVjRHw43QDzofgfe+koIZ3OnULZXIsBA
ViSDRoMfV7IblydiFEBe4WSxvBGYOG6WxGONA+MuWJfFHIeia2O2SUETHYFi8Uzp
eoHp0Xt2JHJFePJfZkCvgzWQJBAHF2umePS6aOH8V3i2qpCSE1GRmjTu0sERkX7Z
GG80ezAscV8Hvvv3URfpSiey7AH3yv+3xPDlRbEgBhJ7jRjlpNl6bmqaDvgCXA+O
VSWx59KLhgrToj+uS7e0v8lSM3zr29C40V1p6idaDtuS9EajYOVMQpRf2DkOB/yz
QhdQUpC3W0JzP5yBZbHwEZhGlmGmKVPX3Y2dVuog3vK2ZizfpFnPh33b7r6/V3ef
+iM8bBD94MRRKwf8ZyU3qzy4iir6hhQbLN5P6K1+JfNkQ66bd6YTdby0H/e2EXjB
Ungt9kobsOZikXnlGH2ZrgSAADN4hNS79qVQgrqdz7I91KAfXsZkrBPVpFD2bUFc
8/t0S0p0kV1BZQ0ZYUC2MY8mZcO+fa2H/8pdX3m0pzm/81cYHyEiyASVcTWCYBQE
kjuM9IJNGBL+BnrlBfGfUKsL53jtBgqe4UbJdnyPhJ9fVyVKIx+HGZi82xeDEzwA
KSsG/wEyWXJ+Jc2bZnz2y8qU0E666TURe4lgn5Hx1fbQXEJOSsjJ17J906FbHXQH
+h5Am4fXyaqH1tztPcw4RcGdSYqEDYeyYFWKRb9qToQjMIg6vXGP9IwHif6LO182
lVQPh4UL/iUA5fZbKwdNkgSMcVJwuhZL1N31Y7fbiZKyEOoTotXFR/GpeuKnEwAN
w+jb8WWR4EBL83aRv7Ad8bpnqa+ZhRu2X9ziKakz05GQVrCqpw3FbXEWTR3MUOb8
TOq/u58OfcEZvAk/sAplcLY9Zwm/ye1r83p6xxewpGHFLlb6cZxXKo+ieuvR+FTS
kKg7UHor+Lev1I1Pt3GCp76xprsRZvVUOrbZFP6GuQAxkhajdMJhGPCjNpZFf8xL
SgmNCPMV1KIHlRTWZBvD+YCxfb+AMDiz2WWAn8hVsWmC9BibUf826qrUAsI99cRa
YUv/WLF7apODlfvges4bJMIzC2LM3RsZqgudy2EhiBRouLbgRup/OjHDxp7iXfst
i8lgoJm5nm3EkG17WP4L5rrpjUspqD7eAp6pRycqoomkfYioKNY0U3B+Cw0dNGmY
9LAot8byPgVAUenSSV/2o1ZwjWXJQ5JngCusE9FOLIuicNx8x7JlsrtPIplttxcT
zfInqxkZBzcL+0AJau0RVyzCaBQQHeb2P/ee9hCYFcnHKyDW7gasmTX2YICFSUo2
i/0qFTLbQ8uf+00knITioMktHJahwTdl1EIvzLEvqEV0STN2Wj6FwyHuynef09ZO
ptUKkhW5IbwjKrr0WS/BHozfNtzgSZw6oRsv4Q1P0ZhXfLk216CMf/b2kJuEsOab
LZCyVUpPm1TXFDhc/TF0sZV0/XHuFBoj+slvtEcWFAlUNjMLIc/6QUSSSlGD4w0Y
YYqdZcb+0Oe1fGTxd+VqaIIfkRls/7RDf2Z56C/oropsd6YYYdLlHZWoTAkbLjVd
m2KUP1Pnt4MLH3g7+jk6GTTI72CmFmZ00bNiXjZEkufqkAOEvZ7es5tUkfUVexVX
6YFDCe/u1K8KWin6KVdif3AwvUdid4jBPzEY0bDBzTQIC9R1j/6a6Hd6Mgrd9Mss
J0u+PiDf+TmxoN6FtJzVmzDk51QzuvrGMyXykxzqWVSVmr63dbVjilhV04tRPqGo
/e5+wd1EmjxO6ZfFNGptHWa7DGOpFn6kiXLqbaGYYhQgNJHEkMXfU6o7BMC8vb20
Ekro7JEHqsRb0JrvofHFadX5e274q1DGnjZIqHs+jLv1LpTqo2HclcWojuCInVeU
PyxrhOfhg5z9WHjlovsq0l0nBvPj6wPhhLvtNj9u7/qK+4NhVoYAE0fgeoNIourn
toSEertImMKkITdaT8JubxbvUicQq0sP3fBBAeAnHAg/fbN3TuBOH/qPBNrsI9eb
OQ70FIIFoXrHOcKZUCCGSLDJPRI1xQoO/osKFPiPJuZ+wmyIi8iNCVJvwQEZe0V0
ZVJnQZ8f66Txp+DvF6hwZdRDtpSUGU7s3xE/JyPJVYYgesb89byUPXfrXEUNwal8
hym20sdUP0n9lyEGuJrGCg1LXg/vZT0XfJ4Wmczp5qR3319Oe3NdepLNl3AstO4F
JDHbehdWQmUS15Tvxi07vbgzpRo39mxy+5UmU/oDh26KdcBnoh0e9m9s03tPGVK7
c0BpfkwwhcWYLePB0gWoXrlSqUSLwkhr8L/v5ONxeeRu6pJxgzmCMOQN+bbkY+cA
4u5jDWGOH4X5sZZRTFfptz3oxFQJgJprhJpo5lrQMIR1OGpsh/MEoGk4ieGFcyRT
JndXRNy6nzRgBWRY3qhWh/wpb/+d5XZNy77JvJP67JPX3KKuT/tjfnVZXc71ONZG
gkIBLAGVfGFyeuaSXBCbW1DAFw8DAExoM1LSNP3et33boC710KfRyWIpqkdCPfVR
DQP1BNmD9DsSZSThqKKDiC/FCoU2smQsRf3DlXwLg4CUylDFDgNta2Mj0bIN+gXo
GFSatPWBpVFHTxdYe3m//jFSE6Unw1ZXFs2kqJZqPRW73nsCo1wQqjUudMXhQYML
RGpLTWxvzul6aNbEIQQPqc+4HzSp63mmkxydz9i7ewhW88PeFhOWJEGYV0CAKMRn
u3rciqw2m5C5ewJOvUDEo6bk0HPYtWxd9NT6ATvKDPVVLHF+5IsqMvGcQBk6UUlS
GKfupZWWRo0lhyy9KmsG/453VA/VM1eZyqRrw8T09zlsVgBjhns1jvAhyTBHCNPk
BmxL3SWojHBQNQKRHa3xTNxUUyTR0aWnfnW0wLFr0KtIH8oH/6eaBnfkyH8USQTJ
673iL4pGQhXHDDC07CugFjARzfehVbbc53/ISxduAM+tjedvKiBzK+aVzrBzw1q2
gFsC0ZMnNgw52i0yGTgRB0/gM8S3h2vF6uYdLQs1PuaG8qUCE+OE4VuE6NrCIxwr
DyFCLtEMDsBQxtUFl4zICrt7UdYB3LARf2UZpOJiivxxcfy3CiuRzuOgdHFOxEwN
4sMVPs+w1pZOgwfBnBtv7rmK3Ijc/xLMfjng7YMThF3aUYL9yhgJqp4q588XprCN
1YTBVsOr7JBSs1i9xt+ym/RiOGRDFtjVcgdxdtovlP+SYvQFnai68/QvBHVM8BEf
zIF5+ZWKQ+eiXNkbj3Bph3gi/KcsW0ZkerRSvxAUkFGfS8egEKH12X1AhJIYAq/R
i7TOLFGuNiCZLhmC80peiaUmEyY5X0QqH1bdRgTUF7dHyTZfAuBAWJdVXMy9sH0u
wYATmC3/kN7r+oIU79O7ysF2DCisx8v9EECj/BykQJkEini0wTNZSe15vq9uu9nM
oxoqU+hlJH01i8JCMXj2doheF6TtK+8uG0R3hMCekUHER8QSFL0hLC6muvGXunHI
isn9HF3aFi1Hy00nKOdervwtP4U2MeuOHv5H4PDHO47E6x+HoG487QE7ajYyLDPk
EF1FX+niILNEk7bC9I0e41IqmzBih8rrDDG9NCvFSh69zAyEbPSQ2AjVW76H+qqL
QlTwBryqry0Gp5RrxoY0S3Ea4GiboOJ4HB+sX6J20OJ1MRFgsHfAkbFXMrw5iB4c
8+0bO2az4xH4WfjsY8OXKC4OSBydd3h0iEiax9LYmDMhktp2YGF3pG5DlQSiyNFX
NsR0hwiYGOM7ieJ5d2d61AzWWfOINyh+kyUlfUKfVRZ7hMHAobuZ4W+OfiZ093By
fh0Ugq0FdxRD57aVhjl5AS2fag/Z+0NDp6MH+rihPsbwL76dNBdTEzQYsYN827Yc
LNDoh8zHHbUdwnFW9tmLt9+IAGQBVt5c0aYMNkJXMQMwyrzSHaQKomorxMmyoZfH
/Usp2kzCKIx/VbP7LeFHzcaAZEI2RLOALyKh4ESr/Gs8lx/+u9o5UNZ7pyITTEOS
2kvfuYdVqaWvYZjvvsuXHi60lVv08D6IHqhM3UW3fRNSuThy/7mwo0h1jqC/q2kF
txHlIRlrCwNWCyd/b7aDjqrgTfbtHzavtaBj47tEk3CNyKz2/UBt0zu7nGQon3y4
0uF973w+96RFlGCOadQ7Ov2/GTGSdvJ8pOtHZI8dYNxRfsIqttxlIfj6ki6uSMna
bl7wol+DMZfFC9kp6ah9m4d0DxamTiwmDZn6kCKc9YQI015SVO65/hJb5swEqhoD
Gm1KmODezn8DjlUR7KsQu7pOkrVBSONu/Eb9YrKU/5kFBJOKT1MkBTqrP1JsHlFN
TGwUQCc6VHstOLRVrBv64FVjgI/DrRfkOc+mLqjm6U2sM8fMMp/FQv/fHbo6Yeui
Aq+wNBW0s+YDNPu9sNr2odS+xJRS3vQ2flvrsWlsy31bKmu6dC8s7M8MHPjmg0dr
ELEkcMb+TXC30RNpsme5yvZCtTI5qpBOHu2jrGtODmCqcFSW7BW6ym/GZY3XLGdB
3VkncY58ixkVJpIwCifaa7uOSx2RSrFl8zLDDK6zeRN+92nn7W8EJZpCwOKWgFLz
3PD0zKK9bJ40q0b2S5HLnYDAWYDvuk65qC97ufq2acB0QSa+akCyX4YqhYF7yjyN
+MudzMoL9rum9V8Chv+fdgcktBwYYPdyAJVSZ8DOVBpvOnLi3Sn/nfhaxBrPy8bB
vrW7x9pyG/lIbTmxV4EfhspYXKIM+jU9LeG0CeD0VgCVVJKU1/4LIR2QCvDu3aPZ
ZcGuQvkCM1ur/I2oX/dc8mb/5VlFCjSNXZSHl25Sqxo+BhhOpCSe8QP9r+l2Ybte
1xwa46EnTxsQa2mvnLzjdPuhUOFooyg5e9gSAZsBgRvzuOrc5XOsZmUaNfquS7zq
SFuKdjlp4cnqq6V8dkemuAlUe1rnoyThHuqa/UIRZvFmAXG9lglbjHDwSzS/j5/s
Vvf9UjUMryQa9Dz2wmCLABD6HT3XxARTqFLaxgMeLOrE8Z2n6AsqUJ3+t9gXkiGf
G64jk4IwxgmITbQlUc+u1XnH9FtjebNjcJeWy9BoaWXglCHXGdQD++gh4X66Pph+
f8KnIkH64h7BCnRICwVMV6+DzvZKCVYS+Dzk+Y3LUNWFPDI2euUdX2duGVwkdmTy
O4WB9/Ha+1GPTP2RsCEq4lu7XWMifK29OiL9ynzHtwb5mQ8WC+XrmOtDZ8Oe/Laa
V6CDxMgRQN4B6XOSBnC+ngQSQLsTk7k0CToJoWHSui0AZ8t7V7I4Hmlz+zmnFtvH
GjF57xeKtg3oGVQi1//9fG6n61++Kuhr6kpsuhBvl2SeQ/Eq+xW955eDmC8hJFj3
tFcOcQfKedWL/ryAD5uBSW2Pn3+DHZCDFeRKny85LPkV+4jGsQ75c4qRjVCOf80W
9irgUf1FJ1RQahjK8axFylbgeE/YX4SBLbDK4L3KYw5tDC/+b/txcBpJKq+m64XM
XFETIEz6dP9qJYQPMBadMMz13bpBD5IieoNfoGpqB88L4K9XhgCwQ9WdjdfWh3ty
TvMH6ItYnjh54JvLMl+zvrLYNtoI+AwTLnJ63eiLCiRhgQvCFxaE1MYIpjqaGcIZ
QhI0U29Bzs68iS0vTXWxIMGiLvyN3mwb0282koCQ27l8pavtXNdF6D3RNQJCZJlx
x1DBX/fqd4xEjFKXgb94BkYkT9BcEaMTuBrRC21QE4SztargbHCAk3eMx98iGDEF
vT+ccfyewUcaVmtHhrtkFSm5t5xmUlwG2QPQyq2x85bl5wK5xS/XcKdX0x5Iezns
J4egqc1l0LIwSPRB2yypW9uezs9CNFU4YzaKYKcvhRi+DkDdnv5FnRDj63j2akzn
G8447hCL/8HE9sqkQZxJq4iMhWOwgopvdcXUdi5Db4kVYbcIztzKEGr6U4kKBcfM
iCyRWeR4twjpiTsOF64ag+2yj4i5ulXfy179UHU2BtEmG3zv9lpiWB1yVRfm3dyA
1JCDOgwFhckAvMeOwEj7loh/bOOBcwlbHJFDBBP8wUapFkRkwr3db8yjum+/pLp3
Jm9QeLSOLwiZog5vGK8IEwm9+EBf260LChzWYBY10YG38egTcoeLwtlcVfqZxOnn
KrPhfo4CRsZ17EQlyVUmcvbMgRV5Epq1of1ohMgqLp3ZbvxRgeR8zXp7xMfeFzoi
gBy6gkak8dZdSZBcxXMT1wQ/qWRI7XuAbcDgyA4hvtUdH0xCTEG7IajQdaBACffW
caTmI4VfaWVCqXjWbT7uDX6zhXorF1QsAF4H3Y5pX8Whl61cRS5VZ0QEJsU2w9sg
+KNa5iz48kX/OD9ANZvJVgYP5AE63JzRqWTMgYm+m7cz4YFdO83IxcPAXnde9F6w
8RKwVDMmaVWctQzAuNpDkwqAXKXdeQU01HvaPlXUb69ktuYTVUoUW94bbf5marlD
UrWGoWO/qi9Y1T848D4nYEueBg7Z9SBIZbsJeALbCVj8BfXfE4Law6BlYl0Ewn/S
S68rEHytwJbTN9pTLUeZJDEJw7xmuWe97yyTIMBdhcAyQeo0Oskvy5iv8znpCWXj
rJ0HDrpIlxePJP53Jrj3jpM3BgsvsoFbmd+2o0YgbHHUUyXtS+zrusq/SPYzSHU+
o7u5r/8LXk4nkTnX9Tl1kxCHgGCwdQJEJVRIqEsDoPGx8zn0thy6iDbYHGvq/ZsJ
1mUPsy1AW+FUW9YWbDKfidkW5GV2ohA8W3GE2PsXSdVdQyPur5d5+q5nzi+xZzj3
rO6hYu+R2KA3cNWEBqYIFx10oPI2sVT4RhFREMY5US+S9K4/SXEbeaTn+uhIVPyj
Sh/8Y5vRdkrNFolm7WxxedEsUpz6qj2lvxVaDu8KynvWgvO7a2AIUDVKtnwNc09Y
vOmglv7JI8undIZVRVsE3CPlk6n40Ho1uXSSosKurXTOluzlcDvgMnNXUM3U5hXA
gwmuDTzsYbzbPR3ZeBZ7Qefjvbjypm/esMuhBtoI5WDd+l/f1+4PQZ+T056wRaRI
VRZVHOe6q/SuPAP+5nnY5NXY3yZGR4Auutu25mN1eOzCpsfr3nU6Ham5+i8EBBbT
sgKoaPW00cDJAQoa9NthKG3+/fMtLGWrdRcOLwb2ExrP+kNpuC9BHfqigJAiGOps
dVLJWB+4vNN1vARwFRe1G2uhBSAAneV0kzXjcy7+pGQ8kdSAbEST2//hpHdmnWI5
rkulvKEBUADHwdqJW7g0XpCaFKRu/CeQgIdGklw7Ra5ggPN6dJc+ssXZdUYXdsUu
Eebos5Zxd/yuPDu2clyDyf5+xJHL/1SRkhjCQTomtNtKRF6F8EKMzNGwVnxc+1q1
iE98StvYFnGuZfPsQJACAB3++SjR/2Uy2x1tR8PRNbe9FxACEb2Jz8b2Ob6Vagxt
lV5wQHfYuTfAT65kwJFipJP5I3gWkpu7CojqatwzgnFVTYd9VFWJl4nPWgJOlcrQ
kz6T+wtxS6Pzw4O9scBQakl/aO7nYj6xlA3toHBj8cCRsisfR7vkgvqMwgv16liN
K8RG3Cl3+eTjl7wp2QCQn9ZDbEUILCwrBD3WY//Hj97Xvl+IPBmy/iUb+HxnxFyV
xDEUCOS0dZj+lfg5lv3KOSte6KtDfiATEd4XvgNlGIH9qNcbeEC6nAVPJxZD47oa
eAW5EUxDIqfyEdrR2U4ldGxNrTBfFOXCy0FgfUqfb/x7p2rM8ALdFhT0pRfHobqF
KWjIWz15MVNZ9FwCHzLHkUymbY2ZorbRDFD4udko/AsqglK7xE/uuHVJeHuJhMiD
/jn4LJ9TNAiSQOmfwNC7rewCpRdHqgD6/i9kAbl18rkRpIe0x8ukXSohVLBvNF+x
xmzjbM6uGSWhJMGm3VKsyeUUvX5UuVMTk7IW7J+ukoF4Ic0BtSAf+TKOrfktN4sD
jZocDvqV0r2S+Zy9iucWXlRZJ9B5PGPFljjbEQVRZR5ol9w548yHIeK2elKIDF8z
waeuDbqEYcNt3QmZeUAVb40xFz/KyG0so6bPVxTx2EunyUNCewm1YpA3YX2hu133
odg08W3J1P/c/tPgcJAdZB6/5YoPTY2AQNjjtVF485X0MPJjah7kVjcGt7pwiwb2
0zQRSUOoMrM+Gen8n+ICVeQFc4pSdCDqHsi7yHfajvVg67Mk2bej1BFHFctRR8Ph
/LSBer+JTVQX+o4kKScY7idQ+RPC15du3ugvhgzlRWyIEMAzj8Y65YmY1yXHYDf2
ToI6uK7aumFstO2Hh7SHL8qWrEtDOmeXU1p6Vl8hN/KmlYORS+LPjusTJVWlADaI
54VxCOVHEI1G86HzWYF763UDMDlf0oOP7R9zAGhEtMe6IAUUix38MndNKH579H0N
3S7AqkxUJvfa+vXrDg2gQXHuYZMVS/o5e5CUH1pTrgTg7IOLNOqQu9HqKj0V9yPd
+UJfLOinvg6zCoKaDXx9Q83zHMwyTGFNouIJWbxEH1nwhRcYAAeLlWHVf0F+IPCm
1l0qrT63N/hltSt91k3X9vwkFOxry1ztllqkZWR0oqJ0JAAuUkhTm94X9i2cR9b5
zwdVQGl717WDwnR8I3jLLS64ogVJSOl/yAwt4nMCC8YT8PcvQXH1JmY2/vxTrZkt
YnVb4vdb3AnmNHxNFIvlMqIf3wVIVR9+K/eQy0K+ad75vo/9H83hdn+T7Jfx9x6v
SRRee9Mfte+GfP5Fg8B/cfDyxX1Y7Wrh2k+JRWdH8sGRFPaOvD/uN2Y2Vq3qzdvv
gw5NgHmWza0grVxZFUkmldhcp/tFW0whr9oKhXdilwEBZKjLY5ImmuMxuaTPzU6L
ExmHbHlcFAOyEnJAZxK+KWpDRKl4TRtOQsQeUS6StpcgUHZvDaz/uuJhwgjEbiIf
dUP12AoQBD+T3HwxNoRIlj5x/2GWPMfQoZf4OuDBTgeyE/s0C5WMXTaOfAR6gH3U
Dq0G++Y42tnsptvHdqZOUSwyb2+61XTxyboA749VG8g/oGGeGiyBngMFGUD5RboV
99x5pshODb/8MY3rJMs7h84VatdniDQMq+s2SQJdeohqdQKe2A9+FzYuoub/eBuj
u+moSYmTAmCO9c3TF1Plfl/J5MBZf/gsvMd12UPmkZ2qFLSXUgJryPXXKUVyMI/I
nk0rk9vqbY8qFeICwFItyRVnV3qqK468Dce4NdcsHnoASx7UywZAfKi4PePO52Xs
2ltr7+kyz62qm4mFSQJUwm4s5yGxCostHjokvECzuSgmtRewZFpeQOvAR54Obv5X
yu/Y13GLqgt1jl8HjcF9IBfE6YUQO4x/APjdIrHKzFM9gaGkZzCCPXhslIEsAJt7
ei4E5aLqCfPAk+DepRIzHiuxjmLpZ3iq9M4QHuN8HFax7T+GfqDy2vn9Ed8UtAj8
onydS3QWArnQzyfvBbU3RJneQlpr9iRUzbxdwa/rqA5uXHrsgxF43thM19vG8vKz
slbUP8vDjtmTX92CkpBBv52AJKEW60lmaqWq1dE9tXafXzZI+nrGXBPFbyQEQE8I
DVxx1sRkbBiGvGLMwkTIwH+1kaooqztN0zTxjDYQzL5IJ3GQO4si7sPlGVs/G8Eh
2BTicqFYlq9H7quwNfc+TKA1id+jiME9aAImWScBkTx/dx/PqFHMWyrevXVc0Qq7
JcOZjz0e0pq5glV5sVnFtLGUvoV/+tIz4cWq6hIGhFRf/fIQAr092vyi8bwM+YTd
baYLaP4t6B1SPwp/LBfx54nqdNjdlZUehTSzVczl+CieLP7N6sU/7GoQ+03Vuvn0
7+Afuw0SsgtCg62mc8S8wxVXnvfeeuJMdKxusvCVNFGNK/67EwrV4JhMm+kqecSp
W/XD48U5KHWVgFvofRjRR21uZ6Cu8KvDKctNMvLmWRb+mYYW4LfwhTWEP7U+X3LL
si3NG6FfyBuQXSIKeUSm9Bdj1H+p8s5uWvQoVaaxOhJsE8om//RJX8YwKdw6JDUz
HKEOLsC+EIuoukYmnVUzuAWpFpLsEUor+fOEpY/8mHVTxmna1IEKHrn9V+jwIaZw
gPH3cxIw03rPi8H+kTYAwmWVPYhR8nSfCDTCVRHP2+191eqRIlLgi1gPAUcYuR1s
VN+24FofdS27l4KaoAshtSafxLIkJRRKkUJ71lvfO3tR26S74PIqKo0MBUqaidHT
oKVffqxFZAuzqDLz8GxLA+ZKMVjhmfXLWLCokpWPiqdcplvxDvfZew9su+ENByl3
uzVCTr9j7x+hYhn8oA6l0l8RVe4RKuftChrdqUqHCm3OOp/as/je+eRiD4qQLPO1
2YQ2Iqv57M5bVkZ6k11DgyVMwmb+0BKe6iKeHL67Dsqo7Lh11UdcabG30suX7gF7
H/29h1CTZsYfC9ZekGdhA8+2pYFgZJOdM34fZXuPnUUZDYrazCRxaPGqMQN1S8d8
dZiOPjz2fgHmFKo9MXEIqpB7RY6iNj101da3wGH/8rsJMVnjVlBy75tfORioKWI/
UEdgafZE+5qiCmEG8EsJZuSUy4BCQ1h4HoCz6HeTGJtIAbkKGiTnGVvE7LJ9osLD
qFK2yAipP3WxmeUN6WpI7WI0fIdomXacN4rd3NNqXRqXCLbRHHvgPh9IIkWqjMgY
PGdg39rsCBwLE8ISog+e+CBdHSfunJKVzQbHi2VP3f6Msd34bnliMT2OdUanPdMm
Lk4m79butezY4LqWAG9ushdIarvOeXzZTU5Oo4WUQ5QkgXYQnHTZg5IPWsrKwCeA
G6TvM+oEf35npDU5YrJ+DWecPs3hPAOPkHW0l8ibL7CWCLb+ooSeJffCMnKCmeV+
uUcSn3F5EQ8EPubK4pyfS3ElAbIGZ+xoD1rGzG1u/ykzZxquz13EI6VArZNI7REo
EQXAnlkBS0NdVJIQ5R6JHgs3+MW/ZmSKAjUj3Ah/iu6NxVLNhYlkBnQxA1KQf7EC
CeXGZzXAk42WhUMjultIJJCvX0EeBg6fZXSj3MtBINdj+izatFgJlRY1aWiNGbfA
6m62sQs8TmKH7zx6rXeT6w==
`pragma protect end_protected
