`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="galaxsim"
`pragma protect encrypt_agent_info="https://www.x-epic.com"
`pragma protect key_keyowner="x-epic"
`pragma protect key_keyname="rsa-key1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
wI+T0k64RZDJZd8HdHHsodDyMfCoJgUZBXytupA9hzpW6lsTvq30r8w973TXFI6Y
pdMhwIjy1CzS7bRwF2Fm06pwYMuj4M0eDmQGOItUzi3ulT5eUHrd95ejj7hmv2tX
jwAgFLutTboK1z80pbrecZRTO5cCZo5tBc/93v57JKzGWR6sGA9ltzKOD9PYWjvC
q2ge5fhcVq5ZD7TyUOYotvdNg7+K7XHD37/iVEKsAy96DAyDTDC4vfOBY7cQhKRI
eGDPj19CAbVw4GK8O+xF26Jar2MK7+bc3/nP4j90xtbZiaL8/M7kqiNl5E8qYshR
nZV20Y76WxFRp5LLdIve+g==
`pragma protect key_keyowner="Xilinx"
`pragma protect key_keyname="xilinxt_2019_02"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
GvCGDJJLOnA12k9J2BUP8F9UQxjtLjNsWMmi+QJqedctL0LXlMafMXf20c4hJl0E
c85Hd0oXdGL64G30sxwKaT29ozTLRG84yD36+OLhsibI7idIQWHu0EvA0kX9WeAQ
c2x7eBq2K8Ruxu54xNDVcUPwHmS9XEMeQkZwJPc2aVqJPocf+5QZ46RkpBPQjqmL
u+H7IHp3gyDT5T3modif+FqpC7V2/fwKX+6mEBkkByQPvsqvCdmlQfbX2DwGEBrm
EkX+w86jVk0ZxI6ySy6vhvvNqh9MONP9bFG00Cgi3LECxoi8w1xPLWvTMf0vCUY/
esulaP/vqcT8PZhT/ELbvA==
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`pragma protect key_block
F9rmDCe6wG+iRSkWLEgVzniFB4+W9friiDBgoNjJNTEy3HQIG0t8AdcnYXDXZZ4Y
SESdkvcR2ypq8w2Cq6MxdxDXh5bVhQ1IE9w3OVAruRx66ZjHmM2WyeIP6Oh9xDNB
cDJkrDieBOVuylBV3ChQP3ceqktWRRRLo8Yp2GrexZw=
`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
ACYsORBrob74RkJHcu02ZOeYSZkYIx+1jM1F0UcA8yrYMOhESVaLtkISuJN5NotV
HMtSzJr6T6V3q0MooTN7SrwNPIYxgszUCeMC1djpf5VGMbfP0s8sem7uedwlFAXz
HlInLtC8wrV7AL9TZ55xv1rvcNE9bIL9SD0oPBmWk6JLD1qcg1Kpltl+crn0M3f0
9/5McBLY5PBe7SDn+ZKZ3qJVOlQj0kWwN0nS7hHkq3c0JIe+XA8xuguV8FF8QaVc
PRlzlWz25wWJmaB930OE2MBn2laNFCQiyqN6Y3OcCdLxk4hPdu+ZsR6QzCp+Hx3g
7imIIuktEw5sOSz9G6n3MA==
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP15_1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
d1qJK/c03qRg/buRHtst4B1hoc0WLFCwtHaRjxn63S3xVym3tVwVgEAstSt887Ki
ZR+/UKhdYL+J0vXq7IR6IRu2DziP6dV6LUF/4B66diwEJCThKpJqZFPY6Fp6RSps
oqPyTTBM863iVdbkOsQ8TazlUHXaK/6Jn1RBXy/RnoUNYAWJO2JUKr2pu7Kc8DQC
lkhrTqDo7uo0qJX+yvU82swASSfViFHmCMunG3OmalU+DrlyYPCar0WmrBfgRJlw
AMusmWXMisUefvRBtDZc+iYCQL04d1gCwvTwi9dd13MDR1GE3NBYF3jNu3reVU9Z
P+jnADOcCr4RVDrUTnjRdw==

`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 4624)
`pragma protect data_block
xw+rgNA/c0ala5WZfAjUl4if7MKT20wb0ChrYyWu+BufPS6lMLpzy1OOIZB+SGSA
yUrdfjBwuGf9qlxNFV/uMOza4DqPtvWKXIofAEz673QluXUzkRPMF+BJl1rP8vs3
lfvVZ/JYb1E6ZvU5CJJ7rvWgnpP/qUCQ7hLSRSiwYTHyjYerY7k71JJ3u2RxlHLC
kjZXr2fU5iTZDffsAxrNvvuXwI2ZdD4jFzsmShbqr4erWjh3c2yVTa+t2RoB3q9h
ZRFxIiSQN0Pi3t64RcHdyHb+vF3AyhiYjzdG7X1VDr7xSFyANiLoj2tHveGjOVTu
lLazVBE1/pg5Ts1fF8xjgLHSgD+ovqd1nWEzTKl1vqtKbL5R6mZPA40IgmK6N9/Y
ecGEW9olX8MYLu7zrtpYBoyS4Cr49waxrtdpi6gb1huA6+AGlvCySoQMhtOJU0CS
1Wu45wLxjwgNgwjsBTklZXYfQyzU+ph+CTD46aP12q8QKes0yG2bDUaYXO18TL2L
zyEJ/53EAm2KovHUNg5+lOnZ5d1W4rsOaPnPhs4UaL4echiWJsXXGZ2aYXTCImBr
Z2FUEGR0VqJO9+6kLclWjaoC6c4b1ZUipVvKpxeiH6a1im2yczyqt5/sMNy3YydS
lrA+S6l0EutmokA97KWiPY/Y0QRVcR/9y+Bry+PxW5vlPolVXTxjJhzWgiowL1xo
K64CBcghhvQkuYZOzzHur7FXZ2SJCGcm3HFK8zM9SZzaruqG/pOYMVrkRZYLwbaj
QRpwFOSWSSfbOu4KVu/9EjmgrFni/O41B4JSiMH7s3avWNi6qWLpo7PzAPS7Yi23
PxTHd7kj5YKNj2Rx6nZ+d1OHxSsECIQkB6hSvtysx2dj7ZfACwXqViTL8lqB86i+
Z+lxpwmGRFnKUwdw9vRF8jxv6MDEhw1JhyWR7AkRPCQMUUcHr0knX2YHOJSmS26H
QBJxKvc3m758Xy39LUQQyzaKptTTJh0e4rMXIfDzDSDYTW57ByDvXpyQj7/MjTfI
TslcK135btaLOysNvQ3Mo65yMo77b346ExXoCOR3nPoZhNzRi4nORBmo3SuiHgz4
gkD8bAhAytveFp2TuDKkmjUHEVBnjUacCLZqIqqWgklopKDCPgi16iREvT5C+BQP
b0OfkD9uznezkvAJX5hAspjiYyJN7/F5+6IhzrHujttoaN+AFDD/TXMS5P/Vox+B
R3BGo4wi6eDy+XF4MA/yLek/pg0VDmerSeXEspAso+96yTT4rddK36t6RSCpGRuY
Oq6vvTNhSZBqH5PGh3mvD/QAIa7O5RQA+6YLURPcPcXUuBAff5taR9kPxMKRMIvg
DsSXHzbuo3cHlitLtNqBefJ/1Vv2IEt/DNtJQFukp2Y45OeY6OwL2bEcxeHtdFxi
eJjAI3Jz5j6baRHQcDArOdHpUdx/vr4NtenJlfHQiX6g0vgonXSFKsxHRhcajque
y9SkVzzqPIjysALdk5vywnXARBqHL9GT0MU9vKsHXYlRgohfgEggKfnSAmhVfBvZ
1kO+kO5GR+5kgytOKh/4AHpOWEAYf0lwib8n1qMTyyYdEnk2tjc+k8Jp1zGNbQlb
wgJG+9SFGx0hXD1nCWVYHp7VsbM0SdQfZA/baII0vVmT3UA4lt6Mszkf/nyqSRPc
1hiekxcS3LboFkJLBxJgzJ1xw5A6Qq8VttDU+B7t0hbzgeUcrG1S94bO7mx8cNAx
vsSzPyYYjKUO2SCgMxYvKtVmjFfKIjYC60xn3YQ9vL/KWXWU5H+ZhhBMIFoVj0FP
QuGJCNCY4RnDOwhtBin1y/msgR64CZqkxwYNQF0Cx7COrRmDWAXkL5O+UBQ6axDM
+rYnhv1ockHjXDkSf5+vzhSumsMb8PiTB3MtWFv+f0u5fpVS3ocN9nTmndi0hcBj
f5VhgUpIwAUFsuNj4ighgow5D7/1TESYj8UhrkkDKbqWAoYVXIeBU00uaTf9Ekwt
asSpFhgHoRKwgp1lNvXvY7fhMSi56ARltV3PiA57iXQLR6OdxIQwJdm9eXZ+Rtzm
i9zEvKFhp94RTJ6jeDfnS//7cAcEimZwy1C3dpcrToEuXh/+x6Gubz7YNTwIr6cH
IIO6kPo537PF20VKnftnTABeJ7yGWdZRHjbKcGiNnzzKvf14276YTQSgo1+GyJ8F
GJrzZigKt7eEDDV5FWH3L+BO/j3Jhb3boUFXQ5oTcOjrk3x5JeFb/O4RaoOQOAtr
g00mO+4xPwN6H8sUnxIfDDb5t9/AICD5PP/qvvmTZ2asSktqbqCsKe8Jc+g0HpQy
sK4VaoDYdkqXhNbX2b2FHv05WzEE6PFMwCc0IxBdaSe9/bYq3YVN9ldmeJLkDBMY
5cM5/BsBKXZ9lbqo0z3BQPtNweq2cFAm1nxHkXYC6xlM2A7z+Fqo12nRiZA8IVpO
WGkm42RxhVdIQhElqdqPbRC4eCUJchbXkZc7kqVu0mLxfrnkqHAsQZJj7sQO8iSY
H2JwpBAiKvzHiSj8bIPqriBfwYyo3d9s7kMbAnUhbsdfATJ8tSIhQxWwsy9kK7oT
6M6fQZG9m/MT/ZcS+bm68BdQxwzZvnfK0Ozqz1CicSGPf8zzt+ctQFsLnRWEFQvy
RZtU+bUORxmk+wC9knbnKRe/gOIwsOefB3ggqr6v42iNFHMlOgAcIG0Pn6Ry1ePi
vc99VWhnq40xaa2ZdDmEtmUjVnKzF9Pd3S51Sa8RLaALd3uED2gGC6IBYUULT+Cq
BOFTzRJiqblna9p9a9Oc4PHSGUv6R077RksSnd7JEywkUJaCav3TZ5SyDYj8pOcc
Z4N3r5BjJBTWxvH2BQ1E+JzkLYYS9yuyacqNYCjbwvE85gm5djvdl770hFGnIy3u
SoIoYb7V03rYPSTNN6LsQ6PMSSOeRjmrV3qVXrYUPL13R9J4EER6FLjyYpDnpF5H
AwomQ5BMgJFgR1TL2xMGbg7qU1Y3DqpxPR1j1ACmqZLjeCpIPD1U3YMPB32mDsKq
zneBjdvzXYSo6S946MGoXC01OPnAENEutM7lZjd9CrxnVnm48jUqDoQjwaxoXcUk
SXdQyxp9LBkoY3aCLuawmnKlerXhABOYPex+JWnzd1FHrQoTrR1CpRUvKZSsXaGs
U/BsC5y4xZGNh2Ua0ZBiMnZkx8X6Ogi2ctA59pBe8Ev0v8MDr/9YzVOLQ1RPh+TH
+g+0huz2PBXj9fVB5a9seN+yk7arc66iskqMVjxA1CQ69tTDlfSeNLxSrCnMmVJV
+X84Fjo1Kh2RMnW9U3kcC8rSLmNzlYDr7bkazzw+7bQyVIxrYOfV2mj5ERWZcqLU
P+4ngn67vtfXSVdW3ESFNfYFUTTsieHXeHnUhKFiDFVM0cPr9YyhpOt2sjs8ANxy
92egjqYl4KfozmNZsMUPe7P4uwV/EboRCb3klfGx00t1eauerwfQx6fzF5gSJ/Q9
yutmmY/CCtjMihF8uoi+GLdmORruBftSbkGv9tu/1hAI0qopZieDhdZ3ub6GUB+6
TIaxKq5nF9nR4VX9Hml5nUxuI4z//Oz3kR49M8XQHNj4cftiEZjPJPyJHjQPr+RD
ve9wcEuUo9QqNR56PNaKcpDQ6Y1IEfxcEcvMXEnnLg1CF3rYu4WXEAEmlsilkmNj
such3ESR/NJ5+v++6cL5sBT7oh251sqLd+iSHopizsRYOmap8oYxPbj1VwPxev6d
3bitMoU1yJWGP32/qKt9Rkjtin1SnAxRtf90lmSKEZ4wHy+c6QjAL88twgQyWis3
RP8nuijBj5ZoD/ZEzlxcVFEUqlCq3pzFESfJ7N5+NiUwdc18BCIucaQEeguDu2M3
tNhuoZeZSBkav3wF246ibGIkWjb8tx91wEhYeSCo/Tb2yWe1TwegwJDWWA4TdHqP
W0pH+oaR8Jjf2/fC0loYCIuCMqmovvQrCYwRYmdgIVNhKIXDNdVJ0jfMldUkA1E5
z7oxZ4qI2DlImHUCOtiGIdbPSHjl4Y/WRV+fJEqy3VanttO7RiJ3nr5MOeuYa+XX
S1/agckVDcMlXFcWkHI/VjNHPnLbLwIUL3gfexC5G8swEO9R2u/sa842uMUjzSN2
jMP8/ZPIUji8p0WpVr1JtVEp3gF7nkSe7m+s+JEys9ZxnZxCklBFf0GbqsWb3fOh
21jV8wvNdSGCFo5C5QNyxiroGX+oo/4Ju3iCnRlsY5m/Lxqy72Y33h/S0jWenmzg
6qRK4Kq4EGESpg+5jfHe5XxpY+PVEf0hKvXicvtw70bx47/auO3gl8fEWSTZv4gi
vgLmsNfWY9xlKCvJ8aV5njIfsDny+D2MEyjvkksZpMbV5f6TJTKaZClR4ZR9yLpu
f2prYNWVszANlHT+5hatTro6nonPpn3Pi5Jc4ElyBs6vFxTQUXzJK6XU2LZwm34A
WUtS75HaCr2owUY5byYIBW34ItxN76c2cd/KROyQU6RaXcktaFsOAP7/cQdm0Y0b
+VhaBor2MgNvmdsAGbUAOI9PwtGhPFbIOnN6gYRC86bNiYCEsbDOtKY/HK2/JVO6
J4e0dkHBa0pCOTmjFU/5uW8eoDZH1C4IncgjW/aOeFqgAzDqBGvOqKDA2uomq9Wy
IJXn0yAiK7FVemxg6IxSPWbFL3b8Jod3jggBqnjK8/TQ+W0Dqy/WaYUa0GFa8HWD
PuFVRvRMGwqTf5qe+d4hc1X5evDcG1eNPB5hItUcM/stfY5NjHOG/WMjUdSKUJ/j
3erjMTwz2azdoPeOOjZ7JCwM1y1yjx7YPeJEK9VeSY+byAdpn9DMtnbmPTICM7zO
cqdjzh7K7ahd9Wlzj8rX2YHuqcECyPptCYed4h66FBd8aQqCQacAA5JYsYrZsBEu
u+WcqyjEKHF1kWraWfAwt8fbafpe7gdS7++eUrejpkXbEZ7LriWH9+z8/wcd5Suy
KQpdcPE/2uNtLBPAfCizJBDyAgRwxC/1NAOffo2rcqEZP9onmcLDyCNyIVA4TdEd
sPCi1dShbG0kQc/69XOaqJITQ9IxElC4BISzj753qO/P8YuYOJvxR3tlSsBwuoy8
Lf0RdRFTDpCr5DGKatM0Rhm5TAyAOCXYk9Co1nO9wDmyr5HZ3rmsbXXFObufEk3V
Gpy+X1BPXKRZ7UxI7s09kkahn69vDilCV7b2NfEdC+/UKqcUF6U7qjxVer334R0Y
LFSo5kuBhGPL5o7fThMhT4sZ7Ul6SHUVZgpInNGLWjL8JJ9FHSuG15ZcZC6oTJqy
5t30PcZNo3BqKJa2twICoPSdTCEILli+xevyNwx1HLGTL0JMf4I0qhAinZIurB5/
DNfWZ0UOgQzb/BdHFchh4qdHHfjnmLY84+2jtc1lpmq0EFJaRVDfSCK8iYWHZck+
/HtXpiRzXkCJGmO7Q+WxjtFlCTJD6lsxb1vmELcNViwLxpxStEnxIhkzWA4AbQXm
uAHN0p/c6Rdxj7RiZvcGMUQbnUdHlsEkaBmK5my9lSvx+BVDTA2cupKpvzXps6Ag
LgaE2Ju2/Ffr7PLJaLfuW84TkdI03W3NM63MgLVpL7+RBX58YIBeojJr0llJidJ/
2OL7QRGc8ZBpfe+Vx5kp65+VPdLUMS2lkHkrGv9NSKLqFsc0ytkl7JZMg6BrlPiY
Y+niDk27tGWK0F6G7uT1F2YxC5MqboXW406DhmEGOm9sOzn0++AkGZm8qjJAfMlN
FQvTZMTGcJH056uRC8WBhvB8/sfBL6Ej3UezULtANJiszflikSF8uW9FDPtUJ6et
dwrewC7RPf6+NP2iNFtXnoLYPxQetl56xwPxfe8F6Fz6+s1GiK8xOc08Lxx4h3Gw
2WvHTcloC8er/aEKHIoW0a7qjIDeh9Z1AYOWNjjc+JblEXH0Ect9AL9DJOUzx9Vc
nQo40kR/oyCEx4Ya20WnuUZ/+w99hWs5ET+czpkr16kCs89UAhOlzTG+ESWEN0OU
KBKndSFiF7sYRIcAoxiVuyCr9ArdktcUt2qw6p+24RqmObX+rAHLuPVx2hX8zw91
7ucHnQKoAuaF9awQbIMXu8oLtMrT024IE1SEd6jEAm7Ek+pDaurPoO6DMbKjfMVb
J/Db6HrmnWzkDwCJIpf/U/hVPeKh9yWOjcsImLIFLtCTeF2T+/+FltB9KibGbZF7
PQzUAe+0XgGUYG1NPgwROg==
`pragma protect end_protected
