`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="galaxsim"
`pragma protect encrypt_agent_info="https://www.x-epic.com"
`pragma protect key_keyowner="x-epic"
`pragma protect key_keyname="rsa-key1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
DU+XyvHwhqbUmxlQYfaekopBIXx2W8FPR8ataOaz4ppQ8Dcqwhzjx236wSKLpCjN
+Bt8dv0+F8+Nv3cWvv+o+fJbConTGjjXoJPBHZ+hsORW4X2J2ITDkmVKN5RAsOD7
3X5JPTjtr8hYz8vz2hiKA8QYtYHjVr2ftoXS2pu0a1EhfcKNp7FlLpUwPLOvknFB
N/Z8U0cuZ4Bz7oCfOfvRzkHNtb4qJx6C8x/WK1UWNDzxZ3AJSS3ZJ89nKDnIxXrJ
Gw3SCvHCXZjnSminHWlFRGeRX3oDXn+DLX9Pcn5nRm9By2tR8aQ+xAtSiZtSsUAC
Y6hhjyTJ6K7lSEgNE18MLw==
`pragma protect key_keyowner="Xilinx"
`pragma protect key_keyname="xilinxt_2019_02"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
OWMngpAyaa3glCOZDAik683xZwZstBNg5VdZurFLKib9CK33u+1MNLconxN9cNFF
b19KFugMM11PiZwDnHcCcsN7+hzqBrqR0dWdMxLzXTH51p5hP1whVlVtVwbPbPgn
sNk7GmKB3uW6X1Mq6+Qwo/d7wNZpRRuQoiNeYFoAfYv4lwksk7bKTnpj3N+WIKup
sYeS27CvBsBJnQnlS3RM6nfnh5HF8atbhxr19CZLygdthtfg7rEz7BcsF52k/CHj
kVomzd+bSurM+maLW16MHQipT3CBDqEq4G8+aeUYvK6f1+XN2drCXZIP0nizEqkJ
P44JtfqlNQcyei/uFBZBPw==
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`pragma protect key_block
ST0VgaqXkHK06V3MUUssTZYACDA1aXHZOLQoA1oj6vLnhp2mc88x8W1g/ovEtYWC
TjB06JHMNXdK1joPvyIa62gB4DZOEiPF33Hk7M+vscj6mqnnoP6E6p7Y6G+RbZot
iJPDrsKDw8je1PVHLlyEjmNz+W2q+GtKKHaP8+oWsLg=
`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
HbLXT+UL8q9Uy1eQDlGlW5FrXN7zLSM07dXfeCKN30gpfCvJAN1LJCbrn8lLRu/b
+FMNdAzp0yDmvZe7/VSv+R20x3ACCbgH2lxnl3HqmFFpeV0UO9pLUVuKiM8ppFt1
+qftuACIinnx/qBUu36ynULD9Djl/vJ8L3L03Mo7S3LIvmkSNUWg9L9hYc30nbmU
l+8tyTAIVcsWavZat03EVvaSsKgCF7+60mVgKNdIVjyAOl3FP+GMi2JOfznAnvmg
RRhdRo8XcZKuQar1iiLU8oVxWYrHIMRINCS7zCQUsga23ruh8LLn0fvtyji7ZNo1
JTZH8JQhxVPZ3xvHpNvf+w==
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP15_1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
mWq1DL2BzRjNbtLlwhYRUgQxWDbGqmGnygCKYuHB8kxeWnYzM9SRH5kCbgB5oM6L
DZV8xf7+7u0btZpoHDSQVaP4jrq1nuczBQqr6N+Uof9sQnXZr93ZXAiSrHAe3c58
x5VlmOdsrU6/XmDsS1PgmcXxP8krYJHlww0qme+TdJ753TBf5oeYE3qqL9+PUOdO
lJJazaYnWGc293fnGwx5tkYbZjEo41+9F1S8/6lk/cybNRkGOHpuY8TUzcvUw1UL
pQ0JVe1lu7lfoBqHlDJvIeKH2HRkiOoqCyVZ8ogn3B6Vgw63WSSRgolWyYbbc/ay
cExSRSHyaIyzPDQyk4bxiw==

`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 67920)
`pragma protect data_block
Ma602q90A0eP57j0LFJFXSvIZ8N2I10YmWHVCiYyjvhe0wGNTsS6Iwg07nseBij8
wOreJEVEHUKQL1ASjU87XHRG69bqRz3peqiRfChD6Ej3sEgs1j5jZ7b/ShVr/kAG
92Gh2ZYNCvv5C9KVtlg3uW7X6Yk53gNmtSRLWN/kJ/qiwoRfYwm1Ycc5rQSw0nBV
kJ5hTSx8gwxHNp8ZTXYsF6rD864xWMqC+U6hhIIsxwWbF1WyDvAx9bc4Mp1tKpO6
4AMnmrELgcTzjCi1BEQzkocY24jj4gekZIhPlcCJmpfwmE6dKog2q9Dqa8dGfb5X
MkRHrxziWPHbWw7uxKlqcWul8snAmUT4p9Ns2NYvziEF5OhwEqoVTATtK7HvQ0mH
o/8/7ey+UDB6wzqiyN3HcfxxJJW96UN+875v+sijFtZp7GmD3U+gvgHrE+zmJ2Ay
AkUkSG3tx6pc7PDCd0kr8AgrJTMbuxKVi59Hfh4ACtlDTE3myKrYj4dE3R+gn24V
lAR9klsZMnANdZeUBrGnF7nMq1ZJMZfZybBc51rQecFNKMGqDqvRxU5qJ8MC3K8Z
As1S4HspP+QZYrCV37YN5fj+FD6YXYLwd6ggCpMy47FMEhBPreB2Cl05ubAvxtqp
iKYGKURtrcdziAfFm4muWbDVEf6yo3TOFKlYQfu8+B/PkPdHtEW2Iuiyh5fGPgVd
T/jT4NfQilNlMNGTtYcizRQ7NSVdWu2+20ew7IHRuvPwZSHHfOIjgsdMbNgrlW80
D6scSuZs1F42EZ0OytfFIbIp6Lp3S6toa//mUbVWa1a6+uLCM0VwKJaEquRHEVDW
NPjWjaUrICc26Y2/nE5kK4qxx3Gb5Cen5172NqLvW7c1nN/IGSAhRvAa1CbhG7kn
EC36AQndnFx7leaZMxOQ8TiR3JseWeRp/ClkXhKMN0GTrOeMRI27Lvx2CcoZG9RW
g/Xntxyinh458EMPTnGXTU2NWvWE9CP+Rk6iUBDoAEI1cjQ1++nQApLo/cdsStMS
aGxGaH0mc9EGtCKHCLETL6ck5Q+zXyQWhMHC9PpdgqMzVeSzMbDSxfJ1vqfYOu1L
DscaPibMnnFsJwag/IKFsrF3CsBzO4Zbt+6QliTicuGpH4XeWwnJ7QvlLgMu5qxy
8Lu85oWklUg+Qhv+aM8eCB5XU0bnylA+eH9O8gRX/KbguquOhN+x9oDOVz0OE5FO
wRCdSOlY2ZMcPwlWXGQZfXBSemSvqIMYFL4Pr+04w0cddGg5whDgBUbSzfJJVKX5
w0vcgF3nyNlYevAz6Gx1CGyp4LWemvzgJkxE/V1hsyh9JlZze8gK9xVW4SAqfguQ
hj1mpm5FAupf4M5i28QyWt7MeBEnk2EsbZY7V3rgZKX/i/J9hPMiYYnQAUGqgyrZ
6ns+bOQzCfggmHb9yrFdzqBilL2blsO+Q8Dv8Lb2j54L6rzpPs4QSmeVMUhXgkz+
PGPD9UjFR2krxrs4nvr/6kKooeAQPGh2VXtH1quhKQJR4w3y3hboNe4xKafB3HHe
37Y2OHoizt4JovHLF3968fRSUYrBzLivvDNm3djPWRGre4h9o6Sg/u+IkxOxfMhb
N7O5RPjgT+O/giINi9IT26f2r6OQ0Tpvw4Ko5sTwthNno9JsPsTNUomgKhHPI74x
JzT/U8VjFfzVIX5ifnRVTboYPVdonzrFkFs/vWnpziLYyQnN5e8iPLG7nTaILC17
kM6PvCIm1Tb7R6a/jcl7/OQj9mjV5/cofdbBXi0FZevguKmMD33CJMFxgCFpsXaS
/1J2Xr9xVkZrOYY/ajOYprOWXzrTUQHTfrwHk2KpX7J4GIiy5eWx0615R6bRdQ40
rex5mh1NoduZxWj6JxTGhgYEsSn2cFj2MsWYz3xUWvTzHrB06oTcfZMaJ3GxDpFr
WVEdl7kVmz3tHa3ofmDAdnboS1Rtj3O1ZYp95vjJ7ogfBMqDFhpIxbRUKp14bcva
Z266Zbyv6Qg6Bq82zKOTookh/w6/XJGEMyKkeuhnDw9N3lAXyafgM/b2woexhTjW
a8QEXCN1vbd9H6qYsXS+4pUHgKX8OLHfU1XEI8L/9t0StOV6L+qC5cJH9sb3qez6
dNUrUGk7lHHje+M4mOqNMyjSLDMAqypBvgj+h2FxPzIHAqXNK2nyJRNMlEJStH80
cLZoQyMxjqM7V3K3+DKxV4mn7UJ+ybvQoICDIaLIWL7TZ1pOEpfH2hhDHnQKeFMh
lox2GFnSX/u43UzMp3sx2hURdRDalripyM8fcPgoQsrHTu9MGzlpbwxJYnIaReHr
zEU7fQJ+RH9BZWoglCuu8vPjtBnqGppj0q2OXDNqbMMYSz+zDknppVcCkgk9Bruu
oFNVrPQr3Edsci27U0IlpDuiJcjhdKv3kUBwnhoPrjNTeGZeuRmQHjvWx6DFyR8z
U/siCs8/W3mFU8GgOfhd4/ft6Bq5tq/xOUguwRtPma/yQsvPg9roq44nfMt53Zz7
PwkKflcgSohOs2G3nKeOnmpg8MQQfDIGpb23YUjH2jAMX2DEj0KU1WDPMIAqSTQR
S+ugkpAZct3ARXbC42/uIXA5TNVhsYoCox0tZ2fZJiBs5iquWXzH9CD0aI1U7iMW
EbkKPY61ruU43FzGQ2HRL+y76nwi1ln9lyqWeoCHjraDe2O0CO8hgO5szmPUro82
3FWkNYYx6zZJwUT1HKqPykNs1kHmdYVnJi3WrkYBK5O2VxKznukRjDz05z4LDu1z
zE4tkOxbm+30IgeU2lYqBG0nlZHPk/GuHEX3PwQxg/2N9DtAPb/xQNTGAEINaVba
PP4/NJUR2bihCPcZ5ytWbAKgRFnqw//ZG3WgYBVceGCWROYXOX2YaZWoqbAkbElH
MpAN70svGXq225Odez5k9XWcAMGtuJB29LqAGMrek48MadwBIJVZOXddfOm5f1y1
NEi8fMkOHP79eJNyvpe0Ju5dwGLEvWEIMh+1D48QQCtieyURylcB/gdrPv7rI6GX
nGa/zK1+h7y/k2o8xDTinfAKYb+ZILaSFm96c98YYuCqvrtXhPEQBbohohp/EIAf
0J4XUvOd5fmoM9RRPoUq+9iYWnokA5LT2gbe1jVsi9hhsY4qG+oNQQ1OyY3zhNwf
E8nGM58EfqdldsTEHS6FUiTqUGjpk5UJ/Ur7KoQZqP3fYJQG20DIJnBkmdC4U3UZ
jPt7nJa2wI8axbNyXdZLOYjcGnsZCxXhIMdPagStiCW97BFUWu6qDduVy2S1fZCG
dsnGShxtmAPRTE/rXfxL8WOhtB1f/Vvc1ivRcBnUETOesvMyvkn/KLljHSh7pPnZ
lhMKxvuJTKdOFP48PsKzbFZRNpr2cjg2eKHr3f4W0F5JLWvY6sFD0vpikwHpC/YS
5M8AZ6X7Brt5PEMGGsZL4Ne7KBWvb2FrDZcDHYdIA8BKRU0ysl0FPBD02MDdMYUD
CH7+BuWWf4yjEEXApxnV6A6QIWn2roRWwzIvfbxHJPsF7V/3Gc4F3meQBiJ1wRms
pYDyy0AL2yjd5mnElIEkLSjmNu0vqQcohCBMVyEPv7+/xWGuaWodQYATS4G9ZKBI
gehAs0ql89SucDcg7xqzDzSdHOqRIH0l3Gl4wfx0p0jK75zmPwNhIS5nhJLeBwsY
cAAfQ7sX8cX5gD/5EV8MGSsB/mJclZwpkelgrHojt8pLFSEUWodlrlxwKDPcAwAk
7Mwh6hU6D/zPTrohjKM6yMWXjxtyUKKGHOoWqCvxg2zw1JE/XRb+V4a3ID9RdeIm
p6HZQibH2R51T7GvsJaiVa9mn5WfE9C4/QnlsGDOyv6k91iO+TMArGbuV0vBkQJs
5lndLvcfxyK+BGZjYiPXY9CsynD9cI1HTsbxgwlW7w2w+gwHvK0RroBnf+7g8DKv
+qRGoWNovvCyo6UGOqd1a845M6TtpUvPYujfMXp8Inp75M2toEpv4jZNtIak6GeB
q6ROM0LK1ks0sQq/tNzNZafIBNI1W7b+nh92O4xuy2Tsj+nT55PP/fMEVqDXee6A
g/fYIChFhK9dF7AFeG23yWV7RUliXXLT78DuCbux9ltkuAE8tVJfuwPuPjfwOXOo
xHg7G9SNxpFhZ61q9ocj3YuH4mCESPWCrIrIHWdUpe/PL+cp1zlkIAZQ+mIYaUnt
gPPgKqm+4+LsBOCaLiO+n0EUw6JlEhEQ6sOE7BXdEP5hYyx3IzNGxlyw/v5Roxon
yQP+9cYjEeqzrfAS5XNGYS6vVx1eSnu5EvRWosIxrrVR7vwdX9nJ8YsT8ZyvRGLH
dRbOqzLCQQLsf2bjA+7GvkZNlLf4yIEnawpgRmO4UXL8EbA4nOFVpeZDJPW2tx9z
0kLM2QzvDXuJka9L7tV9jFZm9aO7N2KVfzCVb6gb3X6BRb5r24MV+qBZ5V3Yrzyy
zrClrbXQuv6VZKIB+BTpDKsHj2gUoJKZQLKa5jKmeZpbE9lV4zh1ZtptTatoQZTr
cQXddBPotgcCnEe5nDL2e7wCqOeZtS16YyrAmBsau6yT6NqnB6OuhTElVY0vKuoL
ipUIAnJGRn+1m+eXs/snDdeVDss4cDwQ9z3Xnpap5g6WOYSObkm+4G9Ryrf+0qgy
+qW1TVv0y8OcxvxQ0lrvb6k+TInnFSG4FvFfaJYenMtKITrDY/i0ne6fyNJWz1Ik
sE3HWoKDioTa9PtM143Mb1j6Fixc8+aGBeMMsC9autzAffoZU7ARvZt1InCC4qUg
hMly41wX/lKbQZG+OaOJJZ7JDn6I6WUIsuEq7sKeHQu+ximRIR9NLf94+RqX7Ppi
67YBIBDXkAOw/CorX5XpLHXg0HJkZw+VV2i8q6d+RVt4txxnrVLhDhUCOk43lFw3
D/+2vAx7I6zxheoQvefio7C4Ud46a475V58hrvpTHwRslbRAqDTvb1ByS2StGhqX
CnsO3C2ZNe99Unibfc+xUBXe4qb6nzMrm6r62OV5IEwNWvZW+kEtx57iQxkDGmqe
dTUPQn8bezD9URKrHOfvrch6P2GvXVAeXTd0y3fEb4VKAjcYVoHDWOiFtEXOrK8y
3fHz8NGdeXD1KXvtrtLU95ZTwaY9L3kvEK5JoEsYltGUKHc4I2p13A+gXq2ox2ka
UyfFBgjWbHbw5zOdNlTN4cD2GHP2Xt/sB4VAO3DiKqfJvNU2190FYDdRUS9Uw69n
E1UE8KMyVyZStebHsy1MerY/sRSWx2P10Eao7Hm0qOWmhFJg7bUtYAqcxrSPGMLp
Fj7/JHtLnKBUk+IL0kzm65BC8nRiBJaZ3Qt8t5+FXBe7X7ZAQOy3nWAa0TTqx2ZI
1A2QSjJkapWEt0aHSu98JounntF+iSqhcOkgWrcHrIhttjUpkxjO/sFgTTd6nVN3
XrjiFFkBpjsldTe71Jzdg8I94XmgQFYCIaPycwPoY/1qzTGlf/4E6MNOZAJpM9Fr
INsX7jwGGMjOw5aoB1Az2E4ZRKNgLwdUDSWfttCSPfVqhhLmaBWQBH0MznxpLgUA
WbxjzlyIwuZDOaHvuH19Lb0cTJTBeOLmiPRHJoPe0NsnDbIRU7oqAXt7jpZ8e/tg
IJT1FeBCwrnaRGNW0kKDdl1q+Q6rYc/V8toIGmqko5NLpc3nc052m3LzNqYLpiuy
hUaP+02hRJizGs5glZ+E5E2ZBTChEHjJkKfsuzbUrF+yrY17BS1WVClXu+6pTzY8
Rc/Bb1xXoD2vLKiw1RHnvodRWMbv+eHZVbrCQfPmd59iDc8Ko/D8BY6xLEip2ahl
0Ig/loZCedFwTIqghshruCG5ZPguatbt2cqQkl02rWqvJttlcgjkXtf+d6HyHjq5
fH3z+lVohdWYpnEZi7kXr9piFr6t26Vi9wt+PmNxPphMPtELJEFIXmDJ9nIduTRa
NfQs/MA+mmeY5ZlzaS/Uga3mGWCWO085VYiGbFirmVy9aN7gCQe6WL9kpIWOi7fj
AcczVm6m/iC87p8N0QYAkAPQk6alLAUcrTDlUbEWn7IgOFJfoHFlmEiJ+f7IDp/C
5JvCxE4pV4ms2mCNFoxdPH2mcA5AVx/oRVYL8kA0NFlovAUIX3l81Krss8RjzEM3
VnMc5wCvHp0Sd0+h7KwxtmyFGAEZhCJhPZaNm9Cq2yNyqifWhZ7HnMBVNlDHgpQ+
evHTva59NaDlKUno77HbbDLnff466sxtZmXumxrxg3tYbdpKUDi7ScmuXwrdKYLL
BQxFfPZRwQkhNdVK0Facb5o+AnlCgUx9PqirceNykFYOgZ4Ui/pWH/h0fKdJScy2
Txe6nLYB19tQL37ritSNQ+YCgRW4KdQ9Nk8HYr+Bs0ODiHEbkaOG5AI7SyhK1GP1
W8sc0G0fjeklBNxy8o0PfELrhsjtCggRWTfCEi52NnQndSIhIoXVUyTU8IWi1JQY
D9QrFRM7COjd+D69nckkfYmIdIhcQPXwkCYQif5FzJSPlBP2CQDDBpqqMhHXXEbJ
JEYyR110e6POTDEK/+WDRyTlUdCNRKXVOv7OZhiWWRYb5HyWA5DwrZUSXJNiJbKl
8BnTwBbsTamuzVRiFHPvhV3yW9Re04QTqSaZ+kNSQ7NIAMuDd4AYhsxdbmo+KtMG
XyyobEya01J4sHKMBsBJuqzO2jA/3r4PiK5Q3ku4nEEfxSw/pL7PvorNn5upg6vP
w7hWTG+1TZSV79O8azpXtSwfGOkLIKP0oAskULt75qA9SrKnqtanusG/XnaFDK8F
i3XA7HPYacpQbkIHCxogKUdagU1m2po+f+d+3/rdep0glx8iJaA/V46lmmOPvKsZ
r7biYZ3Tdn3bwHOIs7ZvidZ7WUW0LivqWpJOP238YiH2UZle7eXgMJPuGxhLwNGA
aU39WV3VKfC4Lh7vTmuZZpz1j7GhhKWswT/jIZOS9/Vsv9k8LPKQhE/CygaUtNY+
HBvBD+ogrOk14hgSFArAWpdQGyNUQu/sctFZ5CnGmStFEdDs5pXoYGvIlfaAZmv9
KGFLFyrjRq1uOo7qCdbPc3bjocLBha2Z/pO0YCZ5b1vncndtOSBTzhyaBQaS+OmR
kV7BCCDCjG+C5yUZeZKIWLB+ofGIRMWhTl2Csqq5m20pj8E3yOmoh0QTf94dsh+O
qA8TdLpJC7hB6CPD6L3xKkfyEZhAudow8SU/u4qKID/PRL2sjZaxQiXR64gK5KR4
3Ww97blvLdu1XWOxoRt09YaLnlDH/vq/9C2rVY/jYaThuJlpQYqKGWuXelWttudE
5OzEJ2qKSFKKBbai+8IVtAHnONm8N4HbACoL85QsJadqOcI42Se8dJ61g349e4Xe
+CtU7VJaXOiNhbOI4rARrjev78mBt6R0ii1p3cFUltd8yBMgdEzifu/ouAqOmY59
qMUBWvLYGZ9VggHdkyZBYpyZUQQt+JqM18xx6Y7C6sP+xMlTNw1cOQUNun+rpEu4
iqm5Wh3YSetRzR3SNt9AYTWi7+d3cVJ1iEv8EQawD3RByybBA+B/RT1frahHTHrD
Zq8V+N+hqzU8KDR3ladkYC+jd6ugirttLjICeAl+dEXfhaZzTPhYUpGTpD2Sg7S3
DkwyZEdTnveEa7i1HyDRzea7ze2Ne3J+dApHr5nmhox8WCaqYPpW4Pk4Y40v08/L
5vP9sEEFrGQUSCyXFba6d0idYfgbZts3/hb2O8Cp8s3vCmoMTDUYWMpQT1+saaOq
alx/UqwaMCFtbMoVvx5cAWNh+27MPQYfHrDJj8uo+9gzIGVwTbVSMaxT5wR8PBlV
GXvpzGMwmc7ZJHclCZgZc224N98qQF3BeX7QeIvstDZn+s9anKOj0V29O5/BMo4y
ID/Rp6Os50JJUNn+L9o9oxSByvkm0NN94x5ui65oWShe3ls3FVFFoPT5VJ3PWgFQ
Cjw9RVy+wuGNHvVIjcZ9c0T5+m3egjoyL9r/5JHAfzDd8e30cYnPeqrMnmTEHuOB
sQDIioHSWq5G+5yNZyzgDmAC0AmculRv3hsqml/7+kFVIzY+22RkjVQt9hsLLagJ
Isp5o99uTOd/0UboSF3BO9K06C45pokcxwpfi9dTkeLz4ZEYsU7CVa+M2V1qcMaS
anMcTBTWcerAFKkXKZ2p5FLZgOxuN4hpi4DZvjKPdoJIk/jE0gHXA32jsN8QyIyr
31Fgkq0M4ADBNNkQVwaVaNvmJ6cd8jZczP1fl+VmexZ7hmt/1ulwKyQCFWspd4Un
0wRuEGrPMjaEtjFpTEDPXqcm07lHEI3CtpUMxjpPYl8QnHgFDcClypTEWIlfdHB4
V8BGDsgck89fSk/Uv1twQ3Rku2CdxDlgIVTSx5iH2J3HckuxKWjjnp4LNDbm3RGS
/421OKOHRLcaAroWtKOHcoh8bW9k0RF9Q25dokH2gRMN3MAsMaqUQrNRG1G3mxKV
6RR7gm3HqTu4D5Y2xzZ6AZ2qGV4X0QHgD0nMLRMxfklFAdqPv6Rp1Y3j9yKcCR/5
AUGGngljSpkj9MUszhjvWw3Nl8PlBna5zy0ji8cic5A0Kp0CGqYr3krMtuTs0ecn
jMmCCSFZwbH/DXbMV395aNntntboyFjkesXUf1vnmVx0oMVMNr7LgduuCWyfDWhL
W4Q2nYae15A4+6AQrpXn72FMGV32iPoAejMkLjGN695/rJ4eHUDonRTcvfcUpDCW
0aK4tXAQRXjUEGIf9uzTSENn6ZnqdIq2cQ/pIX2Q26e9lL4RfbGPTGzBi4m6anfx
akxMJ2j3gmdDYfNs+cma4Eno/v5tOkFB1M95BYbqGJeO6y+NccKeTZYmb/awfKT6
zwORFL8TcVCZ8ju7Qxj0O0J8MxYjTzKHvByrUraNFyaRaC5uQboQKWaC/B/tLJtN
rKtofxecw2twGvAwKn+mxMnf7klXA2aX/Bo5kHe9y1V5xrIM2vp4NtsDdhesWj/Q
6l7Y99qH3XoPKAuSMNWv0mkrAMs2RiywfJZ1CRCEYesLIzUhUdWNwvrdBAEGk12c
28k0txVTzl3m5hEkWQZbuoyA8CCNhcwnTLRkbEi1w3LKQLjfut4IbhLODrsrqkiI
+R2sq16X0niLLONHcFL90dUl+CKqxspZnveIBelgcws2Gi07L1ST2KcuURArRQwW
M56AZF6afMsKXqWnz0G9aiZpG/EyWutG5F3RKgHSkXTy7DrFyyJ8gFMEFeP8wva0
8EFbHporaOEMvfSoToTUIWOD10E/wU+uaImrkwtdoWxPMAbEljBaM9MY+mZEdqY6
1GORmiJVQk8Q7tbNsxWmCJ6sQ5UhlJ87orZ4YVS0DhXZmnIbO9Cp7c27VLRDPsYA
6exNl1x7pUZCPVjYishLUym2XJzC+1fufV83ASbI+iI9pdeVVqL1ffHTmGxNS0S8
02BPFBdTiTZAlgm9lxCAaawQr55aApk02dBHgAHeG/nUmF1O5IMGlgHGUqX4c299
jDnzX20mxmhYoP2B0o8TX33HBAiiP8M06rtX0726Da1pyfEq1QlzkvDLpnhbIKAk
vzuVxzcuQJavCc8RI7mkbLmY7iy6TD0900FY908DDGqGAnXmVkLGDGZ5oyz0n+Jd
4SMV8wsL1OCUsbxZwzBWE416EaxUCoxgd5HnFm+ioNHOdMwZWVc9jhIYAKwPVxzv
FHmqWuT56UfYzPcNllWSAcGDcK4H1WJ+FCZI8Xk6qy4bsrmwV6mh0yMNu77QWOPW
VRg00qj+m+hmRf97OYGBCOzpyXT0Ner/PanzIjrc3Uryn37yYKICU+P20eE/fz3D
z++2LRdGaA4mhcZiW0uGqA3n/oR4eQfgaomL+HCG43pMv8ieM61F7xDid+/RSn7w
D5qvxX13Quoqg5Q9jjCRrU78bZGpTupO5xnFH2qluUKNewEtDlDmzoF71BK6U0YU
HnZtfrEGHdW03UYnDchLwGpDFigqi9K62qMs65drOddM34tzUNacAp5evzpz2+Wh
nRGRl0j4W4ezL5Cbcut5G0P9xdZoxkgoEMDNjVAv/LK0N51UJhoa/JIFLZCkQdqJ
fJifA+S9He1iGIHPW1ir1ktI7+jmPRUx5nZZjeu3xTnBFP30Wab1CQQuJJ33bT1k
E5VqA2BEV+sDhBpXZZRnQDVVolY3yXlJwlZp9pG2Zzc3WEiaYgY21ozjpqIara9l
SxcaVmhdPe4N8H9eF3rlznF8qNTo0k1AQFnr0HZjlEAXIYcZCEkqvCtTsbTVoQB7
/OJcW5qn2/2dtm+71H1e3/lIeejUSR6qNIkjtVEZhdae4VGC1lv+2IsSaJQQviKC
isqagL6CGBQuoa43cXHpduenpBo+bQaD25avTsSROw54Gr/wzFza9/okye6iaC6N
PjvqovCHt3a4bvTm1YIfZalOuOMtnlNOjGiScFF8uKRUGsTtv0NDoptEFSt3kZ19
Kwvd4t88TiSVdIVCbPpP3953+7QHel0v2fSa0cGBcZPvSCoMCMSpxwZO/6uiJaPy
uW9hv2qKuM6kQgRYQPnJDQPyY00cU6C77okC++pyZ6mdgNDP3XdA7z/UtmJok01E
wsUFFWwgSpRElQuJ13Kn0aHNna7Z4ZfngeaEiMWSINyNsSSGxlc3CYMwwpQwxhJZ
ytW9FI+2Eapwzf8Vxw5f8Q8VxYpoX60FN/KplO0pFP1owu1l3hXt5Lh1Qg2x+IjC
ogq0MaJ+ajbHdNB30Uu1iGYWfVTh/oEugwM9nwumei1PlSSElZ7LrZztoFmWF1pF
27dhRPVkA2vnPmwF2WYlVfQRAz6l8Bw///DVFhRo8202NIKi36ZhGLhk3O8a48js
yFFOmzPh1lP4SjXTDMBn73As5H+w6+CuWWVOhIe0AZqaq1jNmsQShbIYA+oRo5F7
WuDyzIrElx0ly/EuwVLpmBnmjVrVZL5NGWSXLFCjqtJcLXeIuFaw3pMyA+YsdnN8
qARffQDoxuoIuW4heYTYf7JzULj3f1gX79olA4RHWHhOm/OapfwXU9699RZ37sV0
cJ1Sty5qIxQm1buN7JUc+23UfT5T/0ftGuzmWgtM3AO++qBus6bYZdLpRyybz0KS
zQcUHmFicG9MJh13e8G17w8d3sE57Htg5Zbl/A2oV8r/yFzzNenITPFfvRhAtZqo
FVBhT34cv0K/7m1NaazOY65QXI4Geg7kbssMYY6Tc69IcwY3QczuWCJ6vNgB+3LQ
BHo72qIVFJxPYBOCrSp45kEng2s4yAauy0my7LWhX0DdDRONshCcEeWazJqu0ngX
eJT4GWpp9U8b+aUIYEatIJYG6Dn2izEUOyPnyBlyU9QncKG83SybCcC8rDv8r+ng
3L4/WhjFNAzedUXHvE2wfJdBLAl30f3CdKJinROxk/+SMeWYXXYywnBXwZVHKw+B
1NZjwkcSNFzxSHpOiE/vv7z2Uxn+e/T4NWbX+laMnN4e2ePPCKpyNq6Y1nZqA3x0
/bCqTfdTKmh5il5ONJj6EMuJRCkOAjaqTKOyjnv0ZyiCBDIxkrGWiPo9zUmi79yV
YsjOP8QlNlDxKd6XXJRvnoxT9f/Y6ZtnOpTJwybaVsqt/Ybl04AdmPnOLP4oRfT/
HXuu8c+uu12eeTcEYsWam9+MY4I5VZNCJi5TpeQOw1kq+dqOFc9VWVEEdbncjEXm
Cuh28MXkrLnOk4MRDn4dJJblpSf23siaKTGOzrlrnGj4jU40u1HKp0jlH4vYgxyL
I3zfsENbD8n061uYoVdgQeB4UUW1vEVKOYQNC/jVe0OoWs9Zq71XM1BDqiCNNzsS
n6OwBMwFLxygAVWsujmqTZjyRoJa2Z31S4iXrxsYgNlVHlRkAe7qc0Ksbwj7HIEP
25gHHFqumSzY5uGtLAEdfcSCe5x3W31w+00Jl5fTbNQdwRW4RZ1FZJRdbr50M4qd
c2bKZ//FijqtGUO8BIIfsXLvAvppVD0nC97d7RwUIGaL2HTpqBpDtJ/nYeeE7WY+
LoSRWBah00agciSOafmuOgFSWU1O7CcnRhPf6mRQK+3RIvwnFOUJ/q7Q05nN7xOg
OHSwaE556Sv1WHuFt7/mZwwcsTKcu+knyL2MEgzjm5LivkBn5ZBO2qzP62LAtGYR
NXA8yGapBYjwWcF5no2MW09AmQCHW3kzwzvh67WtOEQv/3mois/PinPtkMdTGP8/
0jpJ/ShXThFooEXp4TjUspeeYBwhBplitmXffOvAdl2siu48oQQsmp5GOcByxCP6
Fof9Rj/qQZKUwgNeYTwejal4BrGMP7grau2Mys7hHaqt8/+WYTEXZERSx16iEdjT
M/pS65AY1ppIzkLzGivdwHDs45ZD1TR2DLQ1UXJ6fdt4K28QjgWKcMp7edxDBYl3
Lm+qbyegBQ70FQMi4A4jQVVMO9wQR5zhVlFqN1mLj1Ko8AdhB9exJ0V5gjsiYIfF
+wyuq3bn7Qi2oUX3eP5hU0hAMJWbGpChuQLe8Bq2D/BCK1D8ogfTXOQ7sd/SD2GD
LNCVgCSHHbL+zAe/gJcYJ2nexYwSmXxQUQEA3IbQ29TB1TNlDD9nsLKAgd4rhIuY
AfgaZBiGv3aYvWM7GJeRrsef4LxJW4fGB6+LwgSFiY/cvdx4v+DXi1e98Lxnngh1
SW2rqk/HQWCgY/EkcO8it36uKjqHZnDjyoHPNRzVk9THxVRhax/9Ahb/KvXt1H6S
tJJnHPaQzn69IkVS/GOsPXfN81+9/hs5ljVeXjIwOyyX9yoB9w+qzilS/X9XgZbn
wLNoUaXw751kGgH4KbHPC2x3tS69eZeHvZ33b2jWJsssuPtFMiqppP6fVN+kMlop
8QpbtxPJ98RgUk6HfVH+FOyKJEA7Vtp0lUUGzWkGZhdmQEVGNVAGUBqxVZkFKuqu
2aTK0L07cdeS5r9sSvqvlix+z0//ONzoidp6sVStTPlfNakamlpb++PlP6ptTSBU
NOb1WgvltPYCs9SU0IVuseThL61L6qrV9khLw/dlmi1cQ9d7WX77WjgIkwcJpgxo
/hJKQQ9yEXv8fNwxp9GzGdZILFac4QOeqd1Kjr9FqswFRKjgQOsAAy00vk9ClR8/
nUYJcmuduXXBKitmPBLFojI1CzIOlpoN9NlTuQnqS/xxHcmQZy0N7VbokMHBYbJU
GJAbAMfYVhqmYAwQ1Eo10x/pLWxMQzl0IgyUCEgcrYbYOZQVz23pREq0J1klmKUr
UqNuGCgNPS4ruKCXlCPREM6mWG8/nkFjG8AvPMWsypEhbwuDo46HeBDmX5RvO4Rl
OJegT49KEAqzxEGjBnHLerCW+z9dEXmnlbbkpVU1MsEkWhCkphK+3m0VyfMtoWA0
OlmnVrTA7aTt/pgxt08hDSF+cZQCCqfz4dI2v9ShEX6ZJ/cTToFZc+hns2Cli23z
3Oxa73vjK2ZRKKF5RFgE7ncMZqSWX4C3QhOQvHr8+lhUhcQQ/KCg3Fp8P6K+rJ2Q
e6gw2mK5qHGQ5nhXhiKWxGPLv/MAjmxbx3hbxl0bDIDwJUTshF8U7RkabIRaHKtb
cs7DS765KZGP6ybCKPTUjZ8FiFU80/2b2XHF6YzU6oltNEhRH42c6SGEsIZZ4GVQ
ECvJiJia2mbLMR7IvwoPfC146FIryb2mmbc6SY5kq5ZrRaksPxaMBQToZE1POUUC
Xud1ACopRb1HgcZusClszc/v8xccZP2pCG1DLqRd7RPp7Crc2KwuouUkijPklQBB
QPvACyhtKancSKBawlnXJiXMtFJ6T3E41tFWtmxu8uH80hD5wyiRMKNbtAFF+7kP
9LxAM0K8/1m7EmXR8JLB0Dfk0kLitx0lyuSXEFlKSJtjG1yRpxTzg2CvregDUDHu
D5ajO+SKA3PZejt0XB8DeR8TW5cJWjr0oAjup0sc6jHzRRMhYzUEHnt76BkEVAuR
DC2uwshL/0A8hmwpKEJkij8Vy3dUk4ewd+5elaZI0ysAhjSvZVubog38U3WUrlG8
ZzOwpoONDV1Ji5u2aX9siVe+4Qap6aOa61WHUuSobmc0e7g+GEuKrpuYoWjkRs+m
JndGogMnpmgZMu2mKKJhuQS8vGjlaW/yl/Xot+9vPxIP2MxB1aQ+RiRBcdBA9fSb
JWHcKVSY4sNxTlHuw70LY7MgEFIbw1OYVaiRpFTpYJmD+L3ty0hqW+lT4OR5VywJ
ij2L2v7vCc8ehBv3RbdK2Q+1ha7wlDWIF7WyQQhYsZXVXXdJk5UyFu0l8+vccml1
JSQXKge+y5wQjKQL7pJIFdHA35D2Fh4xXES8CQJeVu9Ib/92x3ShR1BBa33CTQql
CuRYSRrlWdjV5H0EMDTrKhchKgph+xh/7LB7r3p62xvhMtBz+v/3AQ8L6rC7Gl7u
n4YZq/u1esoSD/mXzTfP4xb5hJnNqHMY6D9kvX5yN0pG2sWv1AKJFfYRgORo0E4S
SN5xc2nhNAB1ob1zyuwmC+7eV7sm4AutwivcUuH46QVo/nK6nzX449h2toB88Plj
CxRZGjOi9yl3Z34bgCUvhmWedpdgG5TF6Ov2lDDoC8wq26d5zrqUQlW6H62PB3vC
8ttYzn2mXeZ8XSLeELPUkK1I2qYNpvqBI8O7uDTwVIc7IPQ8rGV/eoZBrZJgDSOq
4UWwmhGsCpa48XvnQ+hy5Cluk1GH0oXCPQYnRTxLiQxyI/0De44BzkhkWe5azf0G
mhQs8QxWOEbxtRZQLyZt9oh7Z6l75k2wX21ph0u/df/Kzj+pd9RUAL+eHIPHOxpV
7PxT+gwF5gZC/3JAjYdu5u+3Imscb7LaB/ANeCpLQqZgUMVJ2Hz/ffIUc+JuB/sh
kWUU8WhW2uFZm1THGTVktYpSNVagU1FyAwv7hayrofG9kQZDTDtc6VncCASe09Ni
LEsljy0di+CTvHQrWaYIXlHaSrRz7ff7qTJF+FNQ5NMFZfpW94Lrn4jCMhARhruV
0TXQ/0tvxJW41tksVIHwXMX31YFCpGVA1BmI1gJPC/e07XUQiLFApDJLmJHmnKYq
iXFV/yyNfk7fsTa+/O5KZYADhHMLJF7QDNFqzQPI4k/UMdwqfGSCdYaAvITCXQe4
W1ckU1kHwBXi6A1Ciuna+HoIejHs/jtzLrV6hgpxk7+GunNlA06+cRrEcTbrRxxz
4NZNyFWlDro3hKv9r2vWu9a4RNPxD2t/v/qTQLRvqyXoOktCJCUbow+9FS4AlQ/h
LXcWsynyvRJFBE0FKPrP+Zu5Swi6lqCXqE2e8PPR+Wv73xQV8IBqD4k3bBTqKl2s
7p0sPW6c06agNb51JNg/GDvgL/keW22NJffAITneXwVvMZOnNeVCGFWFKqLiB8WU
smGHNhE0zAv63BafrSBelzuzZHIBlY7s+LDAkaBbqQY/JepZN9Rhg5uT9CMtM9VW
KWEID2ds4rlbUo2dNrWddY1i5Xm5F3409BbjCu6M9Liw2wzU06UlxLMul85Hnblq
p7gtzTfCAvWXIf4rj1ABEqBqV1GByWrcSg449XYHMbwk7+Ad9DWrqlPyyvRsrJmt
G9KEH3pUpOv3cMf+JxRyX5drbvWV+/oTfPMR8E0QBJpi9NlvR/rNtvZVUP0X4rOV
Muqpb/LD7b665/Ye00h4Q7z6xjELf+E0V66qvyjbdqZ4qpnhuFKs9QcfPbQCP46s
fSDkYCRYsLkulamUj7xo+9Zr9Br6dwPCsWvvvjQD1CT115dZrv0/Nhn2WmVHBX+Q
7LUv9kBkimoI00ZdIkq46N3dg3gEnisMUAhu+hhlPSzOnr6F+SSI4Vip9963ZbAg
lLzQDkkmW+W2+0Cuf88eXbZGaqftOQPnhV5uGDQny2GGJ6vmB0pjdrsnyfwFD03L
tfAkIGKwK7zdFd1m5pwHe+wNOzUdWHwotdll469tMe1FANKkYTwC849R1ClDxAnj
MeSu+rkRv6Lnms1rA2joqJiup7sXI6rGhxcyh2u9nh/oxs/sVK9Knyw3CT7B27rx
MiiVWpkkR5jgRLO1DhoL9dy2afrEc+ZINDSCr/gCszcJj14KL2XEU6HEMASRYh64
0NTo1crGKJdarKMjPOQgA4Of3IlbjA2ii0rmgjObpePJMRV7zW8y25onlm/NFLza
tLUqWHgiczpTSiMu3AA3cS3/sIWFGMPtmgjgU3WLTFINTnqu9ygOR0WMcRyFCHO3
Sd1/npcho6YU9mNZyafb3op5VdIU7N56Mh3pQ4rPhrm8x16JyF9XJisk4afv8e6W
TILF+3iQQUtYGgeLIpEYcYtmdlhdv0RtEyC7rZErB0Z8g02Xf+NOGIsh+BkJIxl8
mIBA9WdRH/0suVQXTuVNyjOCqjaujrfRQfenIGQGQtqUo322DDHhlO8cTqf7lD5A
NBlO7Mxrn0c9xwI2AAWS9fEZAtZ1tr4vC1l6mi4FYCaUpvbkg8f2mW3+6ZC+Fv6a
izU2/U8ibLBLnB03uhQvjccj1FmjWP3pIe/5X+x91X6iixQGtId5AD7lxno3rnrF
2Kt48u0jmIHMXIcXR96m70zpSZem87Lz8LYJzeu0A5z2bH5DFzrMlbDBgeVk3MKo
9NGuDTmoZcIHDqm0wCc6/ZxGepVASYrJQKHQihfUwv4AcFhtA0OZRjDs0klPynFQ
ZVB5Trsm8GH488BRhLTAG0MobWXVPEY9w//1WHtNJsNoDlUAhwsX8x+PlpJbH0Yh
zX17bnQq09EJUZNKWf36Yz/pA+c05mR7W8jyZqYwcejz49vEdRs3imLmCnGvEiP+
1VMTVdD+hu9Lz30FKPALRWSN0oRYS4qD3cUy7C/KUEwYmj38R41+5cpdjzgd+SHl
XQ6yIqZ1D3uGC1q86KWo/7uH0viecales/wDT/tBLeg8p1sGGC5ObNih++7iGCEv
OYeGgbI4DkfXUqrwQL0Br9S4P5Iuvn4IZMR+Bxggc0v29/ACq+sdr50HPJW6Zx99
zLgd2wOda+UnzRFxKpKkdzngKbuLNzsPRJVlkM5DMhzX0S7yW1eSpF9wyzhnpypx
SaJkOOFfUrlO6DgKvcveNoMs1QP5X98ZqO1jyfeIBZwIg0C0LSnmomF39vj3vRUB
ZstdDaFfRxaheoXlPOuqiITcEVNQUvCQUm1pX8bEREYhl+xH1EkyM3RT4cjGRyFp
ANWCMGl/artl9Nzw3rBiKvJHAFcooL+r6Bo4Sozd+PDyLHcCtdVPezh6D2H2gCYu
dBChReU4oeYThHHcdP+aHrrh0DrhDFCDDaggPcCgQyhFj+atI/9PuwFANy3kuHGy
8a2R8eD78aGruBtlefuNW2M1ONS/D9oVZhKFXCDMFCRglp1jrgGsfFrHd/iMe+hx
nS3EMJxGHLq2lyDbt2Bw11pJ66+q7EIMwPQk279bdxMltL0zoY7+05fl1UTsTsJT
U689iq913U15Um/zAlxujraUVZyvJ/n8hhDgx3qkxxLQx2ore8gJ8/zowSsCOI5r
j8xQYyomqzZK5zBh+g1WeYql4Zy822Jo9K/bJXWJjuey2q8n3xCIxUuxRoGxk64D
kLpCBXLJn3unAly/XE7NEw2Irx4y3fBLUi8EJ8LaghJbgAMF9cP1eZDBQO6rDvTP
/bktSvtrE5XXFcoaJTDQUloaxSrSiItAFwzjNlyYJT1PBIk5L7Suhb0JPrVtxWlS
ZiTCF8W9xxLDphh226AIW5/Txslu/6GA32HRtZgleA2JPYyuo9TAF//a2EEf2cmO
ukNA1keVlyUbOOgJRTztfjazIlsmAO5MZbwpMB/x9rVoTMqEUIhgVeM0aw0Ihc8Q
3D4U0MmkS1bevxGPa1kS+QG2EksWPOOz7Cn0ktZigWtGsGObBEkAj4oDbT5qGa20
BUVpKvxYiSEX4p5Gqt9PRsR8wWfgtCWSFYaeGCfIPps6lmpeodqhqp5DgNIGHV6E
+EU/MnMnvBhqvwN87ab3KxN5yM7yQqBrIvsHGQGgD8DaoYuM21E90CsgTqj46saY
IkqOyKaP1HdCmMwBSRRiIDManWTHzFwhBkg0V9AzRYrf54nj+aZuUi7YL3MTAfVp
tFzEW6h6c3MtxInyHZ6A5JgTgIrq2FuE0nWK0xgiUVnyIxl8sRI98ihYAkmZhCSH
SiJZjTBcXH17mQ+4Y82Gb2jq0vbIOekcXc8sFR5xFmPiprZx1C8cPTerkaxJmiG+
+4NrCuq/Cvf6SeTccAubm/80ofbh9uhNxkYGmoQEsyVNGwkKnzUjXYei+fhUhAgq
XuRkcaOx3qz/x4AvU7N0RxDCDn+5+xU8AOsm5kVshaFO5eigkLZzp8kkOE8/gwju
bX9YtRC/3konY3Ck2vo/G7x5eCPhu++KUZaEhutSn17pJ8GmiYp2FNBXuPCV5C/x
Ka9s5OIh1wMjeKIpVbE0B5qn1nNIrIqZ/joDjjNrwinUeR9DedLUTgSMLsq4U/PV
N5gRNpl4+nQmBBIyFNf8E6weIu3+Rc8bNQcN4hEGZuDPhh05OSU+6PfzhrOIiWDR
JOc+fhNBwa3OgRMsgIdhprvAMsifidnbqp4cuFZ8cguxnykNcK3asbvbW2EkUfF8
B4Z3ikIQ1zBXF9TspmTU39YpfYQq04/Hy1irLR4K0AWUtsAlfTN5gdPrzd5Rl29f
De/aiZoazDzM6hwKGs0PVpMxm94rEzkpD0nIV0wslEuQl3l356UZZuIIB3JRUhAR
CQsqLXO6zkB0Y4vHqLCi9qfe2nFiJd/46CzepQIM5j0lh0mea4MHOgPO9lSMktzk
00N4297xwJY/n2ExoxiD8gY8oHLrOoqlXFzlln6UnNw+9NgW9RfdVPCCLsyvDx7P
7GPpYTvsvhfosIzWBoc0/MScRZMp2ZZRiVa+DfbI7nYSaUyInPhN4cu8UrqY3oT1
b/lAf3oG7LlePU9ewEmViU9ItrG5DckPtBD5ai/e7H+1ta/DkT00I77DsOGXD5Gy
iV9Aipu7MTvRuDNNs5WFchQrL0xqlZuTpeWyPF32x/SmMPZAzYve9WRCjQZKTfc6
c2+bA9D27bLDq/pR77xrL76GhoerH4wWlaQ26AggWuKlDDYDwvX8PHA4IkVLk3mo
lHVaVdjdcBZ+nHl2zYxK9Sgsap1PBLCCnw0FHpOPOOBJvMz+VApUyO1N12rVImtk
nFH0tbnT3LG9GjdpfefYK8Y/eps/Opbjs8MGoegYc6qU2aimAkqfnyOj454mcaCK
VDkDnCDiJpTtI5PoDCS7UGv0DAnBYPoe7OyjsscPUo2a0Q6vw2lKADj0aOceNP/t
nXyNR1/HiTBU+qEIQnxjE58S4PIz1NaSI8MfjWAjwh2+z8/IyoLrVRHfWLMyfjDV
mIpcPZT4nozGMJixF8ySNPVWl1FwWv/qSGrA83nVvDbRtgnWQ3kWSy2IqtW46rf3
zFymy5IeHOyh2VKPdmRr3r146L3V1LEZpBZzq0crywqmbbi1/JFj+lXtpPCBQKIA
oF0ahkOMZA8nkQN3dKpgf3OYVj86xCySmTIKprs+t9ZKxwmJyOfrcHqIdhTzPxwo
EMbC4SLpcAJ+f+Mlgh2qw8Zj7x2v0XKJRMZZ+OmL7bv7g/CPk6IjjBkXybvvOucE
CIRtnldU2PADsIE7n6qqqfVXKj5JDKxKjy7ui6BpbQopts9w/1t6zcXYHe09YxZ4
WKZIeMkcr3vGYZ9wC60M4nmjaW4eNLiCbqPus7WhjnSZLxcdWPQD2Va6wnnIYxYG
606VZ0n+ZTNwPsTV70H2XhiSe2KwyL70uvsqONSk+ZhwnJ0zKHE9J1p5PoTEVHN/
bYCf1jUoTUZCw75tsE24DlmVrLdXzJzLRe9C//BGaq65xO+PsxC7GSu9RWc2E9oE
4AACL1kn6H2vVmLCKsIjtEKYxzwAEKky63PYtq7CdVoX0A6rUvKTCizNoRbKMFuH
A0YaN/AsZMzzYA4nvXu1lSSYk0Fah5Glvq70lGIPWAZNx6WcYXkSWRP+vkScYlBU
2+JuuSIJLhwFGVqcjKb6vXXtjM/dOr0TDoIJhZjJsJunkWIpwEbKuLWieKt2Q8nD
S0+8gB8X2cL68xEG5BQAKq8a7Cp5mQa05aaw7sB/5lIf+LnIy5/yRubDENRQY873
EA+0OqUPR+FUxmFMesBcryavQzgleSR5m+0vVGqqMKQsthQplUfZ54tN229B2/Yk
EmdwTtKakt/Yd6A/JrgiBArXZpkaAVoI0ejlJyljQ4eC8dbXucTfrqLxdX84A/Z7
4YcaC74Mt72+lQAY8QuT+63DgGalm+6zwaiXzoxOQE+zLvg8UzJGol4zTwJkL9UX
bv6Ulc3oT2mE4NwjE6u07+ir01ILXCZZRKreHmMTrXioAc2nc7WXSQPvuZNl0DcC
KSYH01a//AkRPGUniW6rJwYTtOtbQHyE8Lvh9Bjx2n50xAg+jxQj550RP9RcM8dl
5tNqZeLxJFT5ZycuJHvp2uHth8A1FeSvLuA+gJTUrYVBDFuxj4rsz0mSHSoquOES
MqWyQu3QQCSaHD1dEOSyyQwe5mGAWyCIRAN21OuIxfp0h6vdZTQF7DjuQa2ewbuv
DFiRIAiJL+mEpIdcgQwh6a1XGmACykO/1jvv+hUseyyGo8XqExTi7fyQYvT4crhm
an4l+wdutIhakUG1ogRVRvxeQvHK/M+voU7xbUkUHyabD8vYFcmhqG5ynJ9VqSF+
3cwI1z2zgdpAxtlEtt8qa7gGkS/5MgPG6sYorzt7+05cz+eonrUjPYp++/a2fOlj
7k9FzpE/+nTQL4NZz7g1969mkyQBVb7RI3eMU87VuPqF6nwXWk6zSdtjPbX6bWhB
MOeHgMV4iEkz3EZAd90w38R6/xZUki/dSWGlGvY/kZvz2hhFeSKSYlC151YJ27wz
WUQ8I8DdM9q/hRFgMXETm/Thgm70CUapJa8cu6fmFuFIMAJmh0UBslzBMTiWST+m
BTDSyrEgMDIZycKZfyZEXdAs6KBEqLipFW9C+oGxfQGV34JTu8X17fGEBp8zpf+u
D0gS3e6CKLSw2Q7+VxfZzQkgxBzmLaSP5E84tr96Uva2a/7O3Dls1aXyYfKsRr+k
4ROey5eFTWM3PVPVPlgqqyu0PvODOkEHozEtncygHj4XwBYuXjivLnvTQ2ldOYpm
jxawSugNj1DaKf/1T797csGEDfU+ZXRT4zUJLC1wvuc26qoMKX9ZjPKu+1V0Q8VL
8iFfhJXFgG/XFoxIWVJXnK2Ui5CH1ID+5h4nHGMcmLtDH52jj6D1/0ls0rKzoyEj
7HGEzQi1VfuHhp6RsdCo9X62PHvnoQPyOZZ+enHpeMUKeQvoLP3H299kYaS8a68p
/egqKaqvvov7CPgeSteDlKK0AWkVTsFjBhaBu4B1cIcuAV9rTXh2Kvwiruy8yc2D
gAeEmsPEUM2E6APfwqkKMwA7azAVReBvCzvC6UPqA0VHpZA+CnkzO7/BiWq5Ay5C
+/QNDHh/wF5YPtzUTg0PU9MGtYzk5mmlnHOrIwkU7iu5waQYR2fa1NwVG6iuZGin
zUuFwGLjv22zVi1DWVfZ1v69EbAwHV62D2PEK+VH893WTc/bV/FNqxyFFy7bzYiD
9Op8QQTitJZ31CcUj25Z7rnbxvxBpfITUm3CFR2JloKXMAq/m4UKiA77n3x2Uku0
0+4dtg3bvZJmTxdZ3zQTkscp43Ny0j0PvF/pGu1kU3qcEU4Xn+rYC3kXUbBGO4TZ
r46j9TXrImZqP6ZZXexbx0dGQzXuwaC5LYw1zeIzu5BxO6L0RZcZBXyBxW7+fQPo
5MWM+f2fVqPZjT5epS6jee4Xszxqcy3nqO1fqmoy28xjiyPz3bTH4g0dLAyoHVXG
tsL6KaOk+ZhpzIWx8Suas4elyTxOb20CwARSSLkbBREAqnJ/OuzFxa3uz7lDOSgc
q7wUnIVlBScWKvH4YpD+gjppbxKTUiMG1MJn0YE1mF3Fj/+X0Dfj73S59sTJCxHi
Q1u36N7acXZ8ZV3XsfIwQrLTu3uuSuRn0fycpwFpON7P3feZZypNyKoC/C+TF7+e
u7GqGTOPrbXj9E3eVXQrqKUgY4DRZtVwJW07/RTy5SGOZ2bs4BUKtiVDVmtEVEha
Mcwcr1qAxwDQHFmr4JDAgENaCW8WeLmWred0HxaSENcUB/58U2Y+fJSOxi8BOgUP
xFwqrWJOKth+0QZ2qbTXowOa1r+0Ox0lmauljuy/DCGqGhjiE9WAGuAKiS2I0MwJ
ebJH/+nbTzIrifclZk3aCc/B9uP8/hBCgtAt7miQ0wVRSIPG8OzwHWri9whtxMQG
vnXOM8rg8Vxz49UhMS/dH96Ug2uQ2UygF8a5hc0W6wWECMo/OCLzSAdPmv2rqYWC
lqMTzBVyItQbelYlwaBXbBDuUhhjaXkHR1FgZGxEnQHW716Kt2aBfZ+jycG+ZKwT
OtijemLCe7GViU2NrVcIrIO5hjTpi2rYHKSBd3lOUgXI2QerrwgWO/gjLnHY8Fkb
wSxwZFmAP4z+PyvTDRySFEPshIjm+cNPPmUTp9xNeKhdLvnTJv5i7pLVZ2sFUq38
WNd9d8AR/6P7BFW+RRPI1H+B+zl8bp8g4/OAVRLcSCnLAa0Ys/jZueR+UZP/6WEi
lkJRsi/NGMFXjMlWQ7kc/QPeGO93l9KNc1xb91yfBlpcBdofzbhwSF2QkSkwuboQ
ZvIfSd3sUc7t+6R8s2mSfE0hDbmSyWujgJxdY1x177T02Wu12MMOAHlq1eP1drV8
+f0K84eyQG7Zu0Fy3+SOjq47p8vuTK+56BmreFSPDQ9gPhKMUdZH2G2qJiQCCNwX
slIoOfixybU/H5O/TTQsoKrflHzOGYjPkKIcC0jWq0ucqDa7v034EGC5JzJeJK9K
Dmhny91S+aOD4RbyZ/3NgpYceZz8f5ZJhfGa2J+WpMTBRNOqGuTOeN4sFzKfxpJ+
M+RLH30SBZW30ZVjIw2XMtQDEnbiXU0LNBfxdzpTvIfxDaEoX0MCSd8Y8g4Kfn0v
u3t1UFYNdFeOvPgGSfMCQlEmiUXxJPe3yjrYw5hwadvnnS2muY05vIajw1mwR8Zq
tY24ii2j1LH4Sv4+3LCdArZznLOzICEKCmKZg3iJLGpXVEpAByBcBXNxNIFJcY4f
d76R+DHt0Wz+pDV8HCHE54vQJf+cyQI/Q8384th2f0yc5hjkq461Ipp1di4Huy0+
VSBGe9upeRDOLL/fOtAFhSTFb/TkGwgAiP5AbocovTbqTgTQNf22IWbajnrwsAnq
BahHWOJT88geVS516aojU3A1Kis/PEjFxFcoib7cr3vtCSpSp6rxP6pAeQfBELBW
jXhdTEs4O17kMOtDNGKuSGCNnHz19acUvzu6Vscwf9Oz9UfO6kTIOPUmLxNSAJS7
osuVk8/Qbp3s2pPkTDapYyh44mRKLjl8G88qcauyc5lQYZKJCpzeRa0aledYTvDu
HC31+m3vRVlKiZP+Cwxt+YdI6Qs6YiFaZ5sdWyEHIXqFZ3WHTEj04T7AoncTj3oc
nipyovrNsXAYYBdkSK0kWuRrf17ofSlbGdbHCXqRt6GWElaO276BlFgCA7V3wuwZ
zRsYjusSMAVpyTjvAQHnP9RIF6aumKlOrggM2QfZcWRsytkyWZUepAWgvyMHpS4x
QKbIr8/2cf/3TyS9i94oJmn+vUl9ehfDuMqe8bCCmDMRYu6Qdc+pFF/TeH1PwaHE
Xr+CHeWt5M7v0kF2Jua94vqbd3hKjULobNJn6GlhakkpsLaPTCkxr0RfcecPaNZU
iSP0r2hej/jjvcXRDPuTD/iIeclv/TbGqxZ/sETwveSG0OYA+eIW0k475VUwxkTl
dcd8TOsfOP8ZztM5gA8wAt6Kr4t/oQvNbvbJaQID/0MG5FN5LhEG1f4IVd/SjDjS
5ifAudX9NeEqlyqt8Dv2Yod38aO6rxFIM3p3DhNMs6c+cSmmej/L8Hhn6znLQHwY
HWwKyn2KUJFP0muhn3gTSjrkX8u8iPEu8EV+rmvB9RU+4lMuGsG5eUC5fzVv7wcp
xFVzhUWgWbYgpWZiZ7c67Q6iw4vmfhgxRF0iSRWXUbveDgivwDeDOTeVMDUfqCan
x9UqM+LkPHrQyM3bdQtwOxzE6XoUv93P/3i7j0O2cBe6Ia+X9aoWl8zpW1zQYlie
Wj7MeGhT9dd5Eio4BLRSsYXf8lzNw/7+tuTVlvYadAXmR6X4MQzXwk6mOxRWyJ6w
apyLUqB6bYf1DsZWv/3JmQbmekO/AmrCwtJw/QNsYj2g+uiVQXzhSRqZbSlNSpEU
izJI5I567AJdkmQ6npm/fEGiBZxGj1tqEHCoT12lYGIlb/yrQgVEeS6FS5W491Ho
R6S0NTQLo/YL5CvZI0jOkM97AKjm2rJCVtUmLj474FmfCBDiJJiAalphtBsexHZm
EVwzE3/L0KhCgQj3apNnOIHKuoOOVbL2dfsugQdIjgVaaFE+CI+IiTzZcC12q11O
a/e+Dm7EkEhVEQu54Sj/GYbn1WsuHepnK1awzqsWU5ckTrSHqsIA7rJNIvhXoigW
ssLLnyiaaDJK8ecRyDoR2BoX37DU+T2Jj5lmzbLshUP3gTRRPppB8zjusFGPhHsg
EIQUWgWh/PEWFCkpdINCvnTKjVqWmfvkQecEoh7UXB+jZxTnFN5VwSKjY2ZRLDGG
xJUEJuAxUOHmzILaW/u4AmbkW7/GCXveioL8wnqnxiy5sHu8WJ+rDW6wamkONeKC
b2fh0MvXMunsu162owjm/mOlgzvqCgN1Al1a3n1Az8x+LUWm1cQp91vj33GrYiRC
HubF3eUqkjth4RBXQnFStkeiHFq1heco+VhIwgjdUo+AqyMQ1iZdgprJ83AaWECV
3nfVSY1sqrFAPeOdNbUU0xEzi+ZyzGNj1E6g94BFY34F5WFnUidOIbKq3x6x3Oi5
fbAZPg+Ge0vAVvWVytmWuSjfuNcU/3wOD4htJf71qyBMCR/PYQ8nm6fiz4Fa1b/n
Z20CWZX7+VPiwbzhKMEDaLStvRmZnDbGSSkub7WfMzpGaia+hOW1o/015VfQHGHG
CJ6qlchYmLP5E7ecHU+M5dUORHm9C8fqRbK802x5L3XTRHqx700ubHWz20axzFJd
JZ+4xwDjeW5AIK6gKdaEHMuIGyexQQycb81gwxauiX8VkZcSEkOaDBtQRD9oIPiJ
nvBMvoYP1vhHssCYUdIhOEZxohbu6oMUssP2yr+NVSM/EMCKvKyC+0ESKbxcAdV5
J0NKDgtUjFB4zxusZrWFLYfLpZduw6SLU2kmo24b1c6LVLZOUVplgkQG0koDJtyN
Z2rDvV544l83zoV4KlqOwnp73kfNkNjutok1GZ//GNh8gohNQMkpZK8HFLytw2NK
E8kR7DmTzyoKFK42VlFONJAvaQTLrOi621m38jDuBeZKYb3TA/n2OjIEvblDVY4w
pzXyrtu/FIPIfIkubNzMehb7AMGjMpYYX3Q4cx6w2AYHdPGJYvHxqTWobA5/ppT6
hJJQhjtKwech56crpd0+C3dD9OWQku7T6q0ls6Nd0V3kbaT90LTOj7IlRvBkLQln
v+XiH3Q5SPCAwk6qtr3qKv06kcClSRg+nD8S+SPMQ5YH1denOXckO1rQYlPvAhfO
bEAYeVdmoMGojW8PLUn0JWY+u6ScXX+zinv8w7ovzfvqyay2xisTDJKlpqKegAaV
j+G7fo7GF+GLQQCrCxKPNcMgnsx62XMSdpDKaN5Q8LbNJaCRP/chsmapfAqvc4Or
netygrviRxuvWPIjDTI6+Gt/VDcD2Qfxj+BPXhbfNICOnO2qJjoS+9u6wAP52nvu
AitIPu1ssd5KCBwIyohRYjcE1n1Zu7A+Aq1Ean6rwYRmi7OY4WunaHrzay9IOcHW
295I1WlU+vRxKono1Flv4xSHHWn9tb/UQQttVTIl/X24V/emmBJFUHU+6RTeizm/
WulYbon5KBg2zmn6/z2Fx21i65HeIh1iuGbflzevs0pyATiMa9E961o7vH6xwyy3
Zp705/veEi9xZal8flhEpIhB07pvTta/fI6F3B5ZbGkJZKpcpk2+Xq39tOSRMZ3a
ntTIbud/IMXUW3rEV4ofOVMw2rLSjrd7ygdWpxvyleUjoOEQmz1AqYnOlLCriCon
FDjJy6JgQdUTbm4rQFIIt8Rw0SWvOc4imD3FcHP4uNhK/My7L9gbof4AVrHQJ9Np
0ozrVvVhROxzpn8c/dNpjs1Hm4d9221R1QMTHrtbAa3ZLULJdjPz2ZQsPegL6E4i
+xx/78HEl16qvyMyDjLwkpQvbsTQnDMUYbgh+fuKON6yqCpVPl1Mv8OeZfzMs3An
6JLL51wpbgsnjCZIqMmJBGRRRyIVUiVTN819+UtANDt6Wu1uosbkBHgzAWYKstBl
Roc5uH+XuxCn0FRby4KLar2FsD5eXTeZU+hihA18woUsFWFqpR71YdE1d9RJXtJ9
tJH7Cukrz3gPF2MbIbotjVD7GXHC9P6zlvLlCxTYAbVYoh7VKxWjRj+zUeDknwqd
ay3oPTKQxQ4SQgQUsiaJl2HmfKEzuiNwxqMklj3M0+rS/VioXB2LfhzMm2LdCO2b
xgAXxu7XpIsZ8uBmHI8zfEH5MKcL/xlI94Uz3iHDS6RsmHYeAU+YpJ39UwKzV7zB
KWb5sTFXwSxz3nlBW/PBhLxSyvFSRFFu82nWuV79MCIC7gtWFNE6MF29hIfOvUVn
PrgdslRtRWqiARTtQvNfXB1VOiqvN8HhxM/OjgaCLk9Cwn1QYWdVgROxOt6aUDqo
mhz+vsoPGxgA41MLILeNPXGh8cLgWQpEZIueJ1+iVfxSobxlIhZSLKBvnpfFkK7p
Ksz/qIs6axnrwHciz3TbVUByEQOyZCDfEu6z6dH08N8jyXUXtWXd3qAGLCr9By3H
LAVHu0v/A7B3ZQJuUXuxQHTfCIZC9UZO20IBoTToeOFUrrt1bBzgmiPOoudHNpFm
7AyU2hu3RBfDmYn6CRybDsUj+m2N1BqxisS9PQBB6jB6OInJQIrbxwyh3UrroByI
q3v9/L1xqY4bhBR+rcmDLtb7Cy85T/NJ/z0NmvmPaS3S3YHgUYUMQM8BBl/bdads
4cOX0csLarwO8BZ6ZRXbx2xKJUipGTWaJKpKxMSPtwKo2AW1cT9y7MNaLcveU3bm
FIOal8aBBn/LHQhLBsWwHGSIQDKSETlsDp9rS8Pw1setd0XiGSfheYTI/EZq8qh1
0YpWxA9M+bSt1GICHzWVQgsPA2aqSEFvrLy2PBdlH6fqgrJL95Iy5OfVUsD6wtMe
mowuCtPgiwM7AIwOyFLALqXWAkOeRyLhFA1Ff8bIvbJDLesl1SbveA3kDqmxZQyF
1eaGOLSLWyaaVuZtemKNCmWS6QRZmnRJge+dE2VQ9Wh9qdmY5eaSVwUGheNu8kMC
NgYnQm6t87+YCtsDNQtN0BoNIknNWEF7EAP+b2Fzgbo5CJQ782xabrzMh+b/IM8H
VrX5Ol68C8t6J9owxa9INV5wzNhOYxwvBnAmF2ItL3RBApOj1ggKN18BE08jnZM3
YNJ0nYpAzGPgJ2mPE8TbTYq5ZGu3KeEMg+Vx519ppoXDlVG0irOML8gzEv5JTLl+
vdzFGkRl42yg4Pf0vMcv+93CLDTMCF9r4AgBZ9504KExnYNfnGAQEbRtuxsCSNZO
vJh+sHWx7gMKAnwqLEzcPLGk0FjAdA0Lygty67byXJ413/8/qTl5NCeh4ZdhacbL
+qZKiaed9QGP5wROyNqkyRrx5NY4hUCm+15GZo2U555HBVditS5iISUjupqfWiyd
PVQtspISi80uP6tybH7Mv7Z4qrk4SwryeuhPErGyWmN4flyKXxoPeeXDWNopeqFQ
c1zK3SdEx6ywF/HMBlap92toR1e0kuSbYPNuOcQ4RwBmIenK3QbIl2+ltBr09IoP
etVAzQmbcd3rVhjmClhNJe3+hKblp09PJEt8TZgaH/GICxUxeA3k80EKQ3pbZtZl
DwV82wHmHkX+64Fqs9AOitsiWQzNpF85fn+yoPs/ATtyIUcvtIMfcmyYfYWaldvA
aFvJ4579nokHraJw9iemE3hu6SRatI5/+hiqR13BdGxM8b3lcO74cU/YvuqhwY3K
wnMjo/9VENG9HzRP2YO/Qfu6XnWoFx5/x5ldTKM1b187Zw48AcQ5Hs8HXfLEFhYx
K3okGECFUeoGh3oRmDHYgK7jweVEdIkzIf5nvGUovDxyGF96jB/dKdYvdjxEeNrB
B3RF7TJEjmBi2uDrHdHCWAHm2Q7+h31l9MefmPBwOTVdAIZ78XIxI5YT3H7bKiAw
jSM+fUhp42L4+OmoZ6yMkEVGH6xju115QrU0DApd/Cr9bGgf4HJkhYFmB6xylzPI
8A7qOiwVQssrNX2xCTNnbtMZ+wIoYdFo3HSuCvZYBqOn225B4ZpN48Afr2z+UDOZ
lYoRd81typYfe9/6ZQ01MXBRBqrlu0wUM/58pDiv+oWYqKd/yGAd8CLOZd5bVTsP
GsGuDusSck62KiSsZzR9djvaeJhE5qhnCZIsjjxu4suByGzWd9kTBLI6vE4p157n
h4pHlifwCbE1rEeS1mrT/yuseR8YH3BpXPd1tlwwL2SprEA7YLaUGfUhJHS7VkeB
KVohtRwmQ5+0/QWV++HMT3iFLtHuwWniENXvBLwrAP/bESKxpCGkDLcjNzKX0crp
osm10UYYkWMZgTO4iRnDViGztwMTLIbtNMIyYpMSHAHGpJ7OBDOpXEtMmsglcXbU
wfKA8DEIZEHr9k2ezjJ9wSBdu0bHkLL72Tv0rGzfO7we0O2sN7lkh1J1E7jqcjJI
4eANPfFDn/THohato6FXKh2xf6neT0lhgeI79ft6lLAgHf1nYyLWA05jRXrzFiD8
TyClkz9yK8jUm1+wUmts4Uo6kKvwklc5LaVsPTZ/dP8nvFamtoJcDvExjOqKwv1G
dzgV1o0L55McCsLnYjXzDhl0gzEug5rshzSaoPQEwgWm0Xo7NaA7j6ImPFcvJy1K
UE2wpomz+xwS+GpRtqIjndBic1w4rnD+Au7vUsOHbVC7G5cY3dop/eZ+wKXE8h8z
U5mcw+Z4ypEkXEY5FgID0mQpgR5B5WHJkjBprp01+smdK4m34EVpH5xEpuUIqNWQ
0TpBipnI0iso/o+f6oqIfvTUeCiR35RMGvNLdD+5EapSv+GkbVYKMb9FXJlfUcK7
UouXB0TILBHn3veZnbwEAk99CbL4VHL8XcHqNe0iq22wBYTfofJGpvk0B0Az4Q8R
KKm0T3nX7ztKyhtuYDr+cTPbmMVgyvnHAbdMGUr/yuPITfwaJqRcsdXjUjUK4kbe
bQi6dKw0g3OhpWORaRkKD2IGT14eJ1raa+Er11n59Bfz/hqiAY0EgzFjl87kzpIH
qj9ef9FlJCmDxW3mhb5NYfrrbMexfDZvHrrAxNJwDDp0vFTOeamKe/YpMyLDutHz
tTV6yWg3PUoOuAU1oW9vAqNfpIfnnHrnsRyv4dkvr/LcJPSZXp02EcARHXRknBgC
zjy6fLI9qlp/m+mJv9563cLsZYDcSVfQaMTMsf13itg8+pFUA5MeGM8vg32PKJnU
yZSwIw6VNQlrhOYgRYApSIVd6GB70KRIoqSObJlmikniwACMoCsOe27W66/cQc0W
RN8Uz9Jr9xupwjE+yqLNWeDYKSTWFVo6E/xbFc1ynF1URDwNWsTJgbwva9ZikZd1
ctw8+xQa8PPe1yOr5fgnXLNk5+1D3PxEqz5tQHW31aQc+w2iBqi9FhnQTADskVKH
tac8wdoMejRDOik7mIqn3C0wrwYUiujbcNvSX9uIqYxcTX8EOFxWJJqewdpfRI9l
Fca+gJmnX/eRE8gDW/Ao36+2MM/U4QZRGyAyr77VTPF5e4dfJ6B4aDy6vRMeGlKL
zM3M7wL6aLejtWB6gWlE/qa9lzTFkWjX1E68n1T4KaCoeEPv+0n7d/EGyRy471H4
0Z+FeTdDRwNbbl0qmIcJvXd2ESbJpkYrtVfKRBWNnSw/TVAHzJxz5SkgRr4cd7tj
RGruZw9tWy4NeuIqttS57Xxu1ii1niKYqzezuuT+76hiaHXkUo/7KNd4XBfXrdjh
JRBX5TQwLDxhF4+VkGYdFKX4ucG412orekLi9TJuJ3ays6hlTgo1pybQlF70OyEK
zcQPP203mXnGz71hNKCUaN4sP7FUVdX7mihoIssC2F49nwfBa1E41TbV25wOO/6B
XRjJk6NWVAtH2rYT8WxzzsJE1OCBsJKiba5Syi4hsQ7v+fJbLrHHLeBIHgm1eRkt
XlPyQKK47IfC6rSnwmqAoQbVb0cawx3tRDvRsEpMWUnYkn4JLD28TFwq4LPJkpmV
Ij6XbUr5dbZ8JDlzvFM5nKZDxdUCPr/x/yxEyNLRL3RsUpYt0jJ5EMzqwKpLIuPT
s5b2OygN/WyZNKJt+kbighBRKiryBQcOZDDkgesVX/hxJ1oFtp6G2jmUzTzPHoPV
fMSKZDb8jhZt9RnYfIx2qRMq6YI47cnci5VGiRkwqIvC52FtWlNGCVm78ugqSntu
8OI8dy1GP+fSFVtF97pS5Rz0sOy8edxauKOyQ8ZVjaMEsRhjyQhCMhLJCf5eemjA
215t2FZW+pcHaCTI/k+bfWBQoKW+c5FqkuNwECt5M5B69VZv7GFApZ/b/+yJGxQB
JB2EYzox6nl0Z1MgKFK55lMtPP64aEs9jP5HHhLhhx7fuIr2Dr3lFuwwwu3v8/GJ
5L0s+yyH8c7ILVcm+ABwliP1wnJH5D6qTCmp8GX8k05oznvg9dV8/ApvdpDWBr6k
D47ssHZsAxyJGSKP2jwm17QzJh2Cr65FcpmG4Xngc14v8aSkiXnH9Yns5vcYON3U
BYjwA2M+bABKfNB4CshDs26FWGaZsNTa5Cbxt5fUaOVnhPkCwHCJq8T8I/TCQIEt
OaLFKUtvJhpRo69x3pqanep2wSDb9WPvGH0ZI3Y48+1ZrJTsqlTivnWdGqMI2YpX
7+8cslrBXMaiboFBbYYgoRqk55SSf+f2ba61WF8uAO53TzlcMlOhgqpUjRSzn5bK
9ISBvMKWxkzQRZTn4n74jEhHkQQpOeTkH/1jryIdIfFCEBeEHVS5WbF0FlTD5fCx
lTrUhW+YjOJAWM4G138jAIhy+3Pe6Nyw7CGTUOlaF8Huxq0ViIdDefmmIFYbTLrO
KEriXSx+CakISGD7+b2tOyYgtzXwo89LIoCYPrUJRnMuMOJWBTaTwlV/n7GHrO7E
OxJJYeELP28lFVd3B2QelbvZ5RfqqdE3DnEXdp4q8BMu37c1MzZteasZjNgKdfA4
7dspZINdmiMpRHV8ZbrCWvZ106v2jJkQ4ui3qDOc/fhCNRaNwej7AEGmOusZiPWg
7yc/tvZiEjjb0h/oQPsJZB5OT6Qd3JETfMAM5GcCMDjjUVbyEJm8ZDgOmSb/Vktm
3jPSXnm7UG4yzLuTq1YBRXuXi1R6wMsooy4SZb2jDNq45+zA2mraffN+9D73HNxM
oXOFYyWdzGxgpfGCpt6p/xK0mo9QIYBqL6p/FUsBRwwoQ2hQjsYXjiWhjBjA7Wop
0eXkckvnoE7rTTw3NCoJJJ8EH4dIqVftRO22eq7t061z7UZHnPYCBMO3DXlHIcK/
KV4NvxZ+w5Liv00AGPkwCKJ9IM3rmJ6HZXMvbCm+cntM3Ianoe9WQtKz5wx4VFGN
LvgQVT32tngi7J67eVurFLRk3B4JKTF2LkgTaF37kOxBwouA326qHUL0ndb9KoUW
aSq8uAj8lt5hT6RvfufDXNg55kIeWAeqbIMGMEmzbuCVt1yqNh3o41uVKbXk29wb
tLy5KvX38bqTCAPEvZcjSDRHgT743olj2B/jYTxQve0XBf33T65DSZQop8G9AhFQ
3UVJrzKX0QxCBmSjuIqtHkyPP/dVWOc9dxfkQJdhl3UYJi1c6NOdMSmfyRC49P7J
8tCdMDbWLtAzuKClPMLy6V830CML27DvY5sWmzJMyQBQRjhrnsgh7hMDW25maRpz
DCWRQxWSNJV8KDnDYuSj6ZADXpzyH56uybSZLzBTOX2djqRqII3BuTZElgx0sJc4
QPhMHaeZ810jd1mTkcwaR7DzKurDIIER41cWKhN92/EikGP5Hiv3t/khyiz9p6ba
4luXmVPELczaIZTNXKHf3GYy5IPyZCCRNvsU2Zombgtwc3NtLs8dz4TUdBlxr5t7
Mdv5dcS7qaAQew0BemfeXolH63eWRAgDaUXa0KP4qu5BJe01lwiHE2tAqL7vqK9/
t4PH+oDwWXDI12m21P3ZBG7QQdctn6QV9tY/TX8pkuP3SBSjTs5x0o+q2sVvqEWc
Mqzy1Sn0mCEk8zpRD7uC7xpKb2gfd2M+QcR8ME6mpsyiv1rKyDeHX8kfJ5xzy2bc
8AWEwMAm/EM1Rne2QtZ5nnuCHOb038NT07eCP6mbULWudZZ2QTJ00NHlyLHUlJYL
G8ug0SURzuSnAZtFYICKJRpjAuMKmlv1tEWH0RDqzxvSM/dZQvTYVRzvTBiGStyh
fqP3IxxJ2mKC9IIJQ/diJ7/CK27aLwzVLEZmWPtaP3tHTMefP+Kc3uguvNnXTFfi
TzIuUsH/yp+1e0Ac9q1azTXbsu65SICYAWO8BoRi/wz8q6+51dM3Y3k8f9NcdaL+
vEWrJiwL7rlYP1ZngbTXuYG3GvkqRxunZvOD4TOv6irowKRTD3M2JFrqrLOCj9lc
qgpi0OhYrbVJTfrAnSXSDcj0iD0h+22V27RN+4X7vxMhzueZgxZfdEYPitsjPw/h
2/hhilIH67piRW02DqOqa1lDnI00Jzd0fUqeOGEUmbfRb/GCPEvJZHLrEE56ePIT
J4dRgFuJx0SNe87sGGkwGUbXt2iynAioQyPCYYq2ecg+IL/WAXIJ7t4UyCJU/5El
20+L15Uugn7xJuYr8X47NwrjrELq5zZdIVUWSLqUjrtEthmY0AUtuQ5PP7Kn56rd
keqC70fF7tLAz2cC05rT5zTI+kVvTn81FdpJxDP+aVlGyxhVOWz2Kjoh5FjwpQwv
o3/hAgvBhtUzT29AnASi3WqRyAbY/HR6U3DMPYEW8S5oYbfuwdM4/9WuxT9XmFEM
tT7JqQzagYnk0i+vmke0vCqxaLepdmbY54BlZDAcHqiU4RJ8g/4NNQVfpYcjqv+K
MVeQ4KUIgw7Vh84cqt5Wfv2JxxRwY3H4dhT9TEaUFRpOiow6qyYQKsR9ROBnpHmi
mtEKc6ULMo0PT9lxdbsLbqJ6kseeYuZ2REpM8h/PoottP22QoADiFGP/qt8P2gNl
dB/cSP0JSj//UeA9Ety6qvhK82W3p9n7wl085kHLL7TR/7s6m+W5iP73neRx4j2n
6lBV4Y8Chn0KE1XJl8pRQ8ttPHD4qYQwuOSx+kFQswYTUNVSmFolyjm40C+2QQjk
Kj635vtzfb+1ifjZvlryPh4NRPmDLdp5EAZwHJTMrL0elrGlXsw4QIC8DP+t1zkH
LYfdd4oXTFFr7ogDyZ2ktY78oxtVKyGOCJ+DojutxQm3UE0x09kBkGL95aHJzRoM
uEI7zikCMHLvbvmsJv46FlNWhXrW7kjHEfNn+sb2Pni4fBzblZnnaJupAWBHdqt9
gNLHqzyD/GNE7JS1n+gSG0R+zrOxunEadVYaD9WnAJbTmUr4FUOegy2TRU343dYm
rSKhH7gvV33burIC0PzaxT5P9OtpTumwKOVXUea3nU8ih8XCsIh4PY8+zlUCo2Cb
/MIMYAbuEcky+h6VWAeP/66FTtrFhZ7fTzFt1SnYxquuwtySLY6h9FAc7O19lkV7
jz0PYLeydO5JSKcL8kvMaCt3R9cUgxXFnWnjDTgPHxD00KJt86ZIuVzsYuOAuUvk
VfhhevCfMAVqszglS9J7Ldlp/zvyCO6H/e/LC6xXNod4UX0vC0sUp4ww+1/KiNsM
N44iqyixrUk8VfKQ+Z+H85BuZqMEOuu+nzLxoIBWW+ewLlAdgzPoK29EjBJNvlkH
Y40xQ8yXdJsL3847C2glK+3rguJQEQSHqTEnaJaD7/958ypXTbymjoMjUXtZgLq5
RlfHdxlM4iNxZr2/YpBfu+2X0YeVkep0VzjeajESsU9penwEVzHBbbA4I8gV6+bm
z318gQ0OCg0iEmApM+aUfHGxdjjIxeDBEVTJd8u4+0p+w9y+zE4jJX86Qm3aMuda
w0MBGglfiwNszzvGwoo+/UsM/rutTzSSV/uO5814+49U2tZk5aBHwK0zJK77V4k/
WCYOroyQ+IeoTyeXoloTKCZ9zTmUeR3EfLXAir/y7hwXqQ5cbOhMfV76xQDsPdhH
hiLie3EvyKV+Fae0Zcu6mJ2MIfBPsaTC4c93JUfsBEJ5gwM20/WjBHVGmIv1Snsk
/4wekpVKQzzI0b77gmGJ0F7anV41YujZT7SKQ9G8LND+tDHv00gA7x5mMQ/yxuSZ
hOZfp1Qessue39u3Ik0ZMSmKMQUZpN/L5CdLxXyZK1UR74ioBLfaWpYCTz/aJPkW
4nr8RD3W67Y3GYAqSzcxxvNuNLYssjr2/8t3jw7lWkh5A6mG2kgTF9gRMe16Ckk7
gus6TGWuXlSFjoXh+9FlsRQqWMrS+UAJJGhnuIWVlFmfA9q6OM+R/fePvWMGfXym
kDTPdp+DKV1JlUVaC3xDj109pai0d5JzsoU9+tqRCo38W5tEIjw3RP/aGWiGpbmc
d1ZnZVmqYfG4JmUwSnR/RY+8YYE39rf0pXxFH3vIbw+1wKR+30pcauJp/bHLd8+c
8nNOQKSzSMU8+3scit0Fh+hTkA4BezMNmaZgaZHc1BzwGzw0tJOJBSnz+xcVF/Rj
FJlGodeoTn4/uXJdE2mYPweGADGYBZMvHHO2qNwVQgGedyahSrDmTOPS4pxk9DVd
vaxZPzdcayXNTsooxoNCrO0tX/phKEohD2pd3FMRiSs7/R0qJY8quG8DWCxXAeji
+qrlc1UqqrOLzdkBcBGse3a+ptkYYgHnH4a6ij8PmAljdj7Cb1wbnV690yCm98M1
E+L9BEa8HKUyrd9Tb9JheSjXag3iLHTLI/YJO79nW195mSzsRLUW+EVwwWV93Hco
sUVscfS1RBIQlmXpmaCEFK4fr8Rzcx7sbmKYL6TzOFwp6ZKyXGtgRYHYw2LuVYUC
xnO6FTg5AlmvGSCF+X9x+lRQuQeeBBCO3MN396yYV20ZYAv5dtuwh+V9RbJtzGoJ
RW/vP16yy8kY3Coy0KrIU3SFmHO6qLKlnW4BPmDL77u8MPTcIeNgVoMhz4h1lXNY
DEjcbVFygofr2zuqhczLwtteJYUAvCBMJ9SvRZ74WiV/IxG0pn5pKIba8QEnwqXz
TTj30wB/jLqh9uOPWRYcqTcF+5T/LIdOlBux2WTG1IHvRUIRZIRe+YmV+RaNfQ2b
WZ2Ox5P7KLDrSMd4Ss+SnwxsW+SyGXBsV1rZFuw+QC6tWERN9ZR0RyYdVs/43FQb
FvLYhmQzBADYPpJ72ciP/NIcZdj3ATB35eCGTT2iDYJ+4cz+3fmqdHFdy9sR9aKA
mgiwtMvY5eVfYQzfH/UquuVAjNQzomK0ZiYZ3LDo2jO4zWkA0/Stz19s+l18Ytw5
B4Iz8oxqvDtjbdzXLWS8oXAvwqq8ZWUJCxAeYxn7Q5Mn2n5KVSXuSmXixNBuJagp
6FpGp91y95+Y+1JSCIwaRqnIoR2qvo9xkCaEDmfJoua0kIkmScJl7Crc4jP9+opb
2TfltiKNHDxxolJ4EeoQf5lz4Z399vZX3bR1xWwqUqSuSVY9BYD2uGHAnOOrMaIR
JEr+an8YOHeiT/QZ6mdfBzmE5iev8BgPWNhA3q0WgAQsfqbmu3ndewTtnEvbQ8eM
Wr3gwR0T8jWc/rgirDwhIS4GONnkHW1pOq+m/Y7FZxvvqX8ufOS65es73RKOxNmP
TVJqe0MwlS1CavsIWQ4hIC2qWKo+4twVf75TzHfqOCobjl03fIPYZnbNsliG/yw5
In2gfrflvCHgbSiwFId1b8FRdjMjuFUUA0kTPTnxCLBXha3GLrpN1LYI68/b1hgN
Yq5BEu3tVYSYVoaO24F/1cEVXSn2k8CYylDtWs4IAHA7nM9uoa1T3LZjk/7ogLRK
iJS+lO1NFcjHS81+lVYypXRDIIh0xMR9PgHIGN0MQHDh3oyDsztagdthHh3SF8W+
KfMxGdgOjMZ1F4vVWHSogcgSWrq1KoQJGswm86UIE2pvZ7MIPwRRSa0LHtD7i0cD
MvKz6LD7CENvAxXGp5RvGt7BVgMRC3rSDR/FhtxcQYBP1izlmUUm9WRagrrb/Y6L
XhpKvWrd4Sv48v1yDuA7r0wfVzp+0ORsSYjwR6bTpmfgOrv5s1gm92P0iIKskjW9
XprMBuLtOI5S/U9A+iiEPJ+ozNhptayHMj2esqDGyCnC38VB/IsIJ7P4fvMRnNj0
b/QV5dQ6U8zR8e3ZKyk8/naZOOc4j2J/kELbdC7axCXg8XdgFgwdp6y5xXdWyGXe
7orNIeUpKHXN3MEVQd6H9tlasHBmnwormJUPBZE235bHbMGzNuYtbFZqpMjyNxLh
5VZGLR2buHlr77NdqSdWIngIbQAcsweecQJf2ILc+CEDbLwUfC0iLLmmdW9VaNaJ
1nXRIhDzZEwOblZ6TTn5GmYqIHfYLzSjsRX8M7kPV8TKoumAo4janeu/Lfzd7soZ
CI4Ahc3w8IcXT3VHV8/DIeXR/nYXeG7q7C8m/Xy6hblmH1efRJNGeiUsOUhrifus
i5dMYXLr6IriUX9L9reYiGK4KQzsovkN8ieFYuOCIJcJV67i4RdYdmBilHG/ozhQ
jRCzNQXr8jrkokx417VF991zwH2Ro8G6lN+QCEyXFUwXaD68g5bG6SoQhqCCDhj2
XDQzL1a6SnofBE18Sw7BD06VDv2W4WWwan529yA4KoDlxuc8lwyBHxqVcDb9i8Ii
F0BOFzrpxsoXFt+3r2E4f3wQ7AVKYJVdHIo5Y3K4gUAZtXBJPh9BXXr1SautVMQL
wNdi5xdK+rOIuJtlrgr7xYOIsc2jJkOLJ6SjdNcyqtfzH3tOmb5+lEnDIKduF5Fw
CO96rNikAl3HilQwk/IhAISXud0EcXQ77e5zdlGfiQqEiz/Nrj+stXN7LYyoSH7/
6iP+Ts8NgcZo/SOZY0vxopf2M4FMAvdnmK/+i6rE+1NcFzJNAxygIVglzmxoL/DW
pYbxCPFgxhHM6/L+00HHmR3A9JD5iER095F2s3oe8CmJGignQRbSljvlE2kf1j65
3DddH10bdLQexUnfbxIbYAzJ6f7aVVCoHaxH+7zwADVjp6C7l7Ui+ms1UoaapG1F
Yxob9v8+GJn5JHtmyzIDayBc4sxvYUdpbIjcIbvhl1y8Furpp6W35ao7aKFyDiCE
ulRFUc3XXoeHVcHYyUiw0DVHfE8g8NjJ2VjNNa3nYf47nLqIm3dSFBVkDKFqzXvf
XYP3d6p0HqqoH5ikCkGyE3czaLfzvI+Lk9zxfgwSR9C7Q1bNP7sALlGqxniJDZuT
M+n62X2UfMuYH3+nhhCE87w8KXqxFJ4hYEMpBrOmy9GPwLABfq9z8YjwuTPCS2Yj
0AeXeylMR8iNfKpuk2ov3wO/nTjkp/UzQnMlCPWSxLNk9kSG68Gikr3rIzYI8FbU
SBTZGObJoUqEpj4uKJpSPPjBv1H5xuP4xOQbY8bC2J1LYrkMkHfsmk7mg0Xe7alw
6S6Kd0lAiLGTZsWSw32S2gjEp/7NI51Uuh1V02tzI93cUUzdECcJfD96io9sCJRI
262/LTU5n4MtU6cJCZSZA9Zq4BtvrXrQvZHbaIZejSTnIwCuCWnRpKy8/fTdsHVe
YJSu9eThLxQUksGKP/BlIX7k7ai3gkYOaBxyH3JDxJ4Zll2sd7HFaSzoL6Z+vqf8
kq+HcE2KaGxSF3yeJ2T/str77ZKtp2rxBQV1Lf6178UjmhIt8DYbIrur/Pmh/jXl
3UUoTs3S10WZI9at7dA47nlDt7eOVXJtGE3Aou+WosnX5acY9PhcQzMgbNVVUW1C
qtYevWBp+iURVkuXJsefHsdQAh1siOd5prtGhaph0HDxasNAal0rp4Yz1zquA+pf
UZo3xfBEsVFDDjSj2j+80f74PBzdjDDEgJHalDY7qyZdG/DN+OPvXfdHdjzMyl22
+G2EEaaXefuQAkCDjfOP2xslkz96dDE+yZsX8An/4urioXB8/2ybNbDD5/6ELbzm
Nze2CKOpLMpYdhYoQIbDUTJs+zGhcIvjJJz8bwuPeqqFluJppG1hmRSqayLK3z5v
1gQajeYMOT7/Y8Vy5cMsi/SjgwK30BWKqFbeRwNmV5QxYS/l2YO+Fachb6CPv7K7
IOi16Plnp7o6hhZ00gdeHO0K7yIRzFYr9QP0IRZ2VXFtzuM2UHNGX1YhvLe5GVZK
yIts/HhhWfrl6n9hxzGGgNMIGx4roZWd5tqxjuLph/QhsdVPm0gNj+wSm2sv4H7c
1wn0LO07VJucVHeYJs/U+VOGpWjK/4AqDvtRDxBS01Aw8diPkcnN022X5XzKObGo
JOerxZbKGymeAOdWKWcq/hn0jZzlxTnbAwniFWS4e2+IhLDyrfEp26u6TL1XpCkm
/4LYqgupThjQdVgORo0WgGV4rg+nsl54lm1QP9XRKNh/mNq4eAnJAi+YiLumrxa/
yRJCowFiEzp73b27Ktk5K0R9pMrE1XhNTE0WPE5X9ZKmsflGus4kiaSCuv9DdL1F
RNOWbDSIcI9cbwtPy+msvWujbg60Vyl52SCAua8baI6YiyhYqTWvoGzJaVGE08/H
NGSpFmTzGr4Er9fjY6sGxdi4+ol8NFHW4Xyf1nznHd5S/aRB9Oh9RITGknnXxmLV
GWDdHRP6y6v7+eHTEbpcPEY3QvM7dHwv9Gc1ddwYhLx0tujLT4fFLGeNOkVTlZEo
iDVx54i5GUhXtaH2Ap9g+jMJTC83aqgUsz2q2X09N/KSV9wSUDk+2Sd6j/H7pTVP
ycz2/3crRHP8BZ9Ef/ESUo2RDzVzlLrLM0FAs4FOm7BFCu/QDYiJKkq1OaS6ggBG
P64godmAQYXmkKhSKFQkydQiGXb+9Rt8lId3rVBlZdxq4/heEd85NOsJzmOIkn3L
zDDzwkjep2h8Ao6nltPEQcIyzgOoJ8GLjZqvTnQQ34boHzDO31b1zc3mx/68j0oR
06Q/OCKmXFwzA23p6AygtyStMwSwNowEauZwZUO0C8Rn37fhqIYohMscdwtC49ZP
qRdziuZurSW+jlfFWjDq4LNlxOr0Pa29ml9LVQP98eOvqWOmFaNzopnodTLr14uJ
spZUEigTaQ6dv/fOzATll4qLXC9pISQ7+pvf2HZ9yd5V2n7Cel06y1eSWVXlMdNg
i8QDoFw/wrNnjj0vOEremKxzTWHoUyC8VVt3M+vrd0fxYmlj2g49a6ZDVh09mqLI
oHUDnrHWqema1RzSb1NFcIZ2gaJvS17mPTVrL8gZ80PEnyxoXmorfUlfTjgvjBhz
gxpz82g3KoZzJwVbMyNyXukw+MUCZ8ri18ALclosgNryIiFJ6BI2tRMSoBvThBeh
iBbA7JNSkdpj2GwQnIulAoIXVMAWlFH2shUjk/H6yNnbaWcjCS0ihz0TybMmff2G
txh/o+nzzcnJV3iVhVszmrKI+GdDu+s6D2gHUMR3rupX3NtPxYZExQfKBDUfXV6K
Qx46VxBp/+onyvHerxteqpnpRTmkzj4cBZgtvPfEXUCE4FBsiopv8Sy5bG+IBYvX
rGnU0pSVg3TPG9kIPj8MS0DzEnmGAq7m1YTNgwUSlWFWwDdcsA1dvcoVQonah6jP
0sbOFLp72y3gTzjoLnUGE8XcOtwAw0yFHQRg1P/MmVFOZ8MozTLtJSZj0WtzaoPq
zUZmsHctXdzeAYWWLItWveN/FhMjsX/hRrlUkDigWLH17nVgF87WZHfOvLvvVw5t
+rdaX1dEzSY3ADxzw1AeBugPBKEkSE0aA8j54P9y/SuirwIxe1FlyCHt0RWtj4oj
JYYjRcZ9LzAfKPxoic7h0DXF50wUMCMGxi/XBKuk6VCkAZ9LGPKDkBUYGqHnCnPt
iYaFx2lDpc19QRZE+c5ZaBfeUkK0k5pFJPO+C4xqyx2FohdTwf7wPq+7xeliZV+X
USjNHQbfuk9Tu2ENHCmrxe2q2w4EiIMZvCkCIO766fcWkW6RBlvQss3q2wyFUq7A
3Cm455ToNeDqjQIuVX8qVhoVRqBbDOxyLrtrjuZT1k33rRDyjdPxWiASiXtUXU9j
C9SnUts9KO3YTBBFFRxClp0ahQuctIr9ht+A5abxSIjsULFP/BWvyRFQ0AtjoZ8F
cT6mQSYpzNS2ROqPDG7rz5vOibfXCzI1HCeUsT+rN0DqXJ8c9nR1cs0A2gWfdOA3
W9ztLvB3tMFEM7nRPofvE3m951EExmKrrT6jd+Bwwj/uM8SMB8ilzmHwiuK9ux0b
vMBlv/DhATWFy/18f3726eShrF2Wt9ZrwLP8SZ6VNrTJR71yWnVP/3s9e8uqXDPw
KKkSjA6C459tu9xQgwlqCTY+LADl3qMJvXfO3O0gezvzpN5CF2Pll1x7jaLyXpZy
QerFjFiTecAw/2l4/RZpUzFBt2UweSX0QY5nBTu2EYJclvl6TaxHViPF7Oqa+x3M
NcUZrlShayMxWxhiHo/dnXEwqGSzNcG0UZq1vJolrUIrBjlhqZY4IREGT03AA+EP
Cn/hzm7CpR5wHggcfcxf1fDvw9MDtK5cWJXQEc91wLxRkY3sU8jo08nb/3wmOHw3
Y1Nyy4jODVXZjz0bVTban0mvxRvpnczuMiU/SfDGgzNTreZEIVnSUq/xjtQ0tmZS
PcC8aysLNPs55dTVJTkNDtgUfScfviGRvTRZpmJB9hy4FPFpvpQ4IqiUwWTjitl0
9hB72Nl/ATk0PZFw84R2xNcGyU7Cgii5fvk+Mf7jNHCZnO9eGNvhRwuB1Huo89Sz
zCgJ44lSMzp8ab4j5YwEQUtWF+p+jg5DrmtVEsS6MYCoMsYjU61wm4JBcjx0tsFo
wtMDrYf5tdPkRm9noaHQkI8plI4PfPwGi+oIRgwvblLRp75JBv7Q2PCo8+p5zTSU
TTZJItsBZEB6qWD+49nrOkdC5AggXg8xXSxtJBaeTE3wywacH8BMZ76yWkmp4Rda
FHGE3iPeCrg1X42eGrmbKWxonl68TjpMC7m0pxaqGpK8jcR+q/UhE3ZaduWGke0S
0SqdxRz/3Q0/EmJm/kQ6xYo4L9h/FlTTJ/ChIpSp5JaAfWPF710wZrOSPdPEhfHN
k51gdrjeuzSP76nw+9+Mcok+CT9q1xIDttwkjFasgGAdlHLJ2gRsHLuRETZbrmZk
NT/0QXrhm5l3oK87T83gwIbFYBkch+l14kN8QqcEne4o8C1+8NcFx+fRRsfTdUwZ
6zg9XP8h6igQQLNqZUvz+/rCY63a9UQ2JPLZxuAdPk4ZrJjocIJQdCRH+eH0huHN
s0SyVKiyG7oekFA0fwR3upd+UeG0WKGIx1jiDjZvTsSOzy3/e3y0d9OP8f7qJEZt
uJ4yZgEgZZWhnM5qCY1Fef2fOJ+ARP/1VdNvwKkf46mEkDiv6YUDwaP4MQ0sGIhy
hQxjL97xrkhZCcvSAGHtYSA2nTwQHwoHIQgC0uObPDA2cRq+hCJ2mFmZ8+p5qSgK
jkbWm0lIY3EnxVyhWrfz5lXTRI6mA4PY84DvxPJNgyQDB2It3oDcwWEOyd5FUKZU
r5LkDLQZhZHPmz38XXFO5LT50FzRr9yACwv6nd+djdY5HYldV8iRP7j0fCzr8J3i
q1n6+Las1LH3caSgs1Xv8C9J4eJT0q8ZQZ2kmkTVwiYw5vUzXv5Q+KNQspHa/7jT
Dwn8F/rY0UWzw3DDoEtF4UzTBFlDfTGV9r5mmhHAsmfwWOfKww5vZ3x9cY4YSTli
lTytMpc4OcJRlm8W+dJEKL9iD3mVvO9tHPwovluLhn6R2CDSZ/NypiaXPgZb73MH
C3I7nZH/9v2Ld/USGOZa2BM+p523ISjZb6KabaqNvn43ewWGLsXOMOS4FCbh4Bt2
ynY2RqnkZlHc0l6/qRd2O+7MfJ3vsUV130WGMU2YvqaL7vsFCS2SvLWvVEwDp0/s
TIEXbiPFryCGGgRxx8WFlclK38S2oQFHYsS6cuOzSB+KpaCdu3YP4R94TnwkaPc2
J/e0InqHND4IV2MwEB+tP1u90HiAEUxqiYq4nmEILVlqb+on12VgIxtXp/CI4E/j
YSIQRpQ68KzOrG1UN6oS/Qo3wsZUIAGPwpLXlxTlgzitvEu9Z1zkUWRdZyjuID3r
ngXXy7q4ArcFFqvxcwZTBnXE8tmCfvDxv0VgR4mhTXewY8kRwCt6t3BfopcPPbzM
pKSo1rNrPAVV/Wwma4BCnOt/Qem9cTxQ7+CdyZHCz2sFT74MyWwD/1mPmOxJULlW
sA956F9qsfsQM7NGg2PWzMmqt1Bd99rUW8nHVofi2UjJAGs83fU14jzCGB7ie+sM
liH9RgeCO07+rGG3WlrHlyDnc9kgQvgq8evInii0irfuDf0lIuRujcgIf939Xsz5
q8Ssu67dOHAiQZRjDTu8Yos2PEV4Jy9GQtyku9YreTI2zLXtazrBrA/ktnIg9XKz
Jqj9hfv9VGcSo2k1o/JKeJN1Be+3N/PaGqCrAvvM8Tss5ojguqI8PiKdIBNYlSTi
/te6hjymR/zO6UUB6N0jfAk/cIjkJ8c7Semq6SUkym0dUlniyh1aZhikFKFmJUH7
+Tzl7i6p0Kjt3fsZAWuDIGWP/lZkEc2n3Ck1vHaZ/uDUNvol/j7GhzoiIZLo+fja
vvjJWWlO9BM+Bue1wXAlohd24BsQBtaZYiTHIf8Kk6J+jSuccg4wbneuY3G7skHs
87CIVm7ZdJhv2CPq/jqBuLhGmQ66JoWu5kikHDrAPw73EBEKxbdY16Be96YWxEEb
6dhgJPpq2lOfUgJ6jLFf5+tBH6Ya4CS5wO4AFVWT0dELYgghuX6AwYRPrLY/Yqur
rtpSvfye1y2JJ91zJBlv1+3K4nKvp1yqkiQIHLWKeh82ag/nl2+/j8r6pWqUsI0K
68j1boycY/Ol/xXZkIhKSd11jZbRbPplWK6vFR9TTq8xIdUPy1UKNKr8V9LAJOUU
3IswwDRStZKs+aQ0DPKRbAuC/8+ETWZ0bEHKHKIeZgtVgUVo8ONZqwMAzJQN78Gs
CkOJYet28eixPCm1UYRH0tjWtIA73FM8BEoca2/YqnBNWi+J+lpaxpdrmzhJvsDD
NHER+r7lw2hfpw+RGfpV9jI1xVEhqPLiWP+BcvBEjYDEcYkB5HYG0IJA2VffYVh8
ru1LT2FPlI9dxG3HKH3WteYjNhkTK2xrFZz/w+/2Lbo2CGIyJNVgOTRGa/w/YCb1
kYhfecsjYtWHKHtu1SqsfCD4rzKkuABZVxZKCwISbXS6TVYfpLEiTsLxfsWpD5Qi
W8pZHqIFXyWOE7c48m52iNMFrNs4IBFH4vX0ALSmdgV716fB72TTVNUUDVtIXs4p
na/BrgQXdGyEgDSxnaneoLcafi/fx5dYuFWIUiZP/dQXv7dnEz9ajKFNBKlA5qik
wtLSSMed13v7yPZeORpHkGhKdi1lDBbuM/bahXQWAvfhpf0zpBetDe6sKz3cT7BT
bLtDw8r5PRaFl3swpsA+T/iVvJxm6OFrAcEJSz0K3r+Zsl+Gne4rBWluPFRXdlec
tIUt9a7Vgpy8Lc6WrapodULZgBtJ5a9oYuc8g3mOnGB2lOndPh99UA9MJ+VWcAqG
eNIzfcVyTllIWVA+dfSES6NthZRFhoW8od4WY9DU39csZvRMSfFOowNDOgrG5hb0
6hK9XJPRRdM6EH2FFNAqQ8IVL9W1OSDePVFbcKNlsC1pXWMUpOrGA/7Z7X+HVTgE
x4+x4jQ1PxzDFDUnh9dmar3i8L03sgGLlh1l5+khSpiaDYnSz2Pq+5fCdzpUSZq6
tHQsZxAx9Mfzt4MUXpw3O0YXYB4SSdsFGisPnhWoaDTfIOMI2+8h9ccRY6fRq1Ni
LSRGEtdL81jjbo4CQAkrFqa8eq3FzT+ry1DdJS0yHBXSB2K64RijxMTTmlcl7FhA
Uf2I4lHuHkzK6SwjZVBnEuy0WY46zrzIhCcUrbWJnyYxmOijEWiR9pQwypXgWEvn
GzzOEefaKUL+rp7GZGcXph4R169g5EN1PywJWmXO/EvXERUmHozOW8Xc6+Zf1KiN
Y3MGSn492fyHHkAvs8vUjIYZIyWtJasc+/kMAR5t1WC1ZJGvFuGGYRzRsnWF98Os
zgkxy1HIPdN1k6VdAEudR027/7WB09YQQalv7zdXdwiamkC1MslswlKj1H1zG4Ng
Gf07FK27kLvHUMijsWbpuLIOhmMHBuIlnII+kQQWIObPSv4kmMq6Lzj5ER7yuf3Z
IMRkv2bDb5ALgtaQhy36WZjMpgcX9SEC6qM2mh1RwyO7T1vNHGIb7AqyuPXG/LYm
J0bNHrBr5DHYIcubYyYL1x4U6xOGIlXym7zT+XV5TjMhRYh4SZpUoVMmNFhjNxZZ
AjdoU94jqaZhOviu2CWO10HkfxNCAHX0F91MixYFQNt1++ZS5OtguxWMgtmDfKy6
s72LW3pn+tXp0I+5ZTjF/v+jh/EWewCKDI3omM+bzuPefKUmqFszcdkc/gOfhRPI
FB5qi3ZC8XZb2Nwq7mZpX5fR/Ya/VYnlWp1Kbae931SEACmmHd4+tLTO0wJ92Ql+
p6V4aKPA7YS9zTcZoVkKdB0OwBOHFLsG2wl+GaSHNmeBGHM86P4kHPEaJfIdt1gd
S50lbRQ4xRe4AlG+zrhOJbf9WXF5B+GkTor2uwSyVf4sDWUqoCweH/gHRmGbsqD8
mX+iaY0fbbZVJfbVksTf4Mj/jiYDHFD+LjvdeQLUf7Dxq3hewj0n0w02EUEwmQpb
4aaznmdf3d/WgsejNhi/mG6M0G9yGL2wQZhMJlL/ZbsamflTbVFHyufv0FpsAKSq
RNAYHhb0ioGPdNA1Tm/lD0Im9fRR2kVCNCOStnjIn16wLkK7tkBpsJHIUjOfQcfA
esjG7W3160PH4jTPqP3XaFoziAmXShRFQiiQjuadzzl2d2eFsllpcyFjde+gblFy
NU0Tq3/emusgUTRgxR+5udeyG0ZophAZ7DgUjF2iC/mYMhWefe3jlrmScb62FLsD
egY5scwVO7GGWiwmvgrM6FiROJdeweiIHGxNmMv8NrNX6qIwfxAL31fRqdlOrn3e
GynDHnTzAHR9/xBdnmMul2YTsOnHUlKDXRJ8Z2IUYFSDuVSALbttAHNzGmuo0ovc
H4buH5e/nV0vXTeDSToHO98HzjfZABW3iMEg4CIcQzgUhRMOKX5N1WW/m3AznBbs
y6pQ/fCOiR8BxJDI7i/Xb4SvRcrz/0q0tWhymDqoijY4NtLV+L7xS1cv3v+f+0g0
Hn5lF+dwUCyT4Rzn692VPkB75N0AmZM0lR9cY+kupEOha5jwg4WkDX5W3oYOxg64
z+ilisdq6RyMkmqNrRjWLsN+P0wDvUZo/TmCGkPWX64P62SnfYWDGJtWxjfDnwsR
NA7QD9Gse8vvdNHI/CimWFW9wSNLQw4ACDOSXVXmccbs/dLHz2pCIt1oyUQ0PysQ
uraz/YtuD8Gme8UhGE2EXKlEU/nwClrxFBoOkdus1o1qdccs5gYvJyZr2nyLq2W6
S+QFmjRyaoJEnjWbO09ZI7/OaEP8hy33EgJ3bIJwti5ggULo0w4ddptbDMulPU3L
mVPZHOuet5EVhLy9sh/TMIHBUaEKtUs2hqcYbABBuxtIMyRw6+fK0KmCzl7n6QQv
+NnDTW5xTQkIFw0bFM6k4Cd8pOWpejsQYola9ADDg9sU6lSqvtcakfXWQ0STw0So
poiBwYdiHIpoLIsJ4VfM4or4Cd4rn58KL6T+7aPupIMEOx9xZVJfBzPkiIj5YhIQ
Rvl5gAmnTmVjiZhc6vrny8oZEu/yFrsHG4c7u9tYGytWdoAbQrOYh7TxDZWMc/E5
+TDcmQK74fUXBBQFsNpSK+NhhRoyALmlZlsAxriM+zDUwp0t+EkEPNDmVtcaxZIq
l9vRDRoHmui4AN9CHwisVeW78WJqQgLq1exREgf4T/84LFhE3n3vsys0p+Me5kmE
XCgTVWXhoT6AGpHuZi03a5fYN2LEtZcRUL2RqyksxoF5zaMTIP7fbLtJaNYVhagU
pf1poI4x35h4fndtZR/5bH2+S+ls3k8WZshFxyb3K2zkKZ5Dk9mZvw1E97WcZBtF
YGwmCvjHlkeITrkgOvh3ntMfhMBfCTKuUbjXH7eHoaEDvoLnpaSYGEXTMUgWJaC+
w1n0vLDlNzwfgyflGOkzdTUGFexXUp48mN/SOkJgEJ450P7k9+yUKVrXq/fJ1uma
nFDbJOwZ4CXP8tn+1ix25TB/QCCf46pMS4uqn7plGccICsO6E+2AE7+aUT8S24gE
nlK1ZuLLeC/RaeRvSv9HguF6srTE+0JkbBAt4bZiZU342dJcV81Acu2jjKl8t9bZ
RmS6oE/g0TBsLA605dMgi30K2jL3R1DyL2fYF8UZAlRy6lJ073BCrJd8R6qxKr9V
dN9urrPOduP3TO7Bn+uycuPlWXCz29O5GrhRfthc2LYPFwBkh0tEXwzA0tHKsBmP
92Kv+ttQk9AsTjEnmhlZHMo4r2CwQZkrhXZAgTgdeZxg+ZJQVclmV1M4QbbqNdJS
0GnsQMftRXg/70bmpmpo5fa/m/XPTyefeIsQUWZXQOHUK32zqpwsAYsx9VFyG5/n
Bmi98KLE2rQotJPeAWqiGg/r9m2VygpTEs7JXgzT2KyAtvSyHYRjaV28CbtA3HM2
KyH7a3XdzwrhUEkGv/Wvwe19qOmPoDC9X5jVjOT8ELO8T6yU2yF4d2fmtbeAgUOr
6vihZwQ1XSr+HSQY0pL0Z+hzSEBiRZxtFubcnm28fzgmAPV8s9KIpEFqysQLD1Ja
j25QpGhb7WufkDM4h8dCfFuXRMud5Vfb/qP10Tm0hXY6ZvHCPUOgHKQKaRMG5jBi
uZ1AIPSO+1qnxiQlJ7MR4H+GS529lO33A8yMs42uzgI0GawThWsnE+AJ5RKCyzns
bfDp+q3VUR3C+Xama6PWN0EFxnTCcDRyCrZHOQkp01C8QUKOa94pMyMXF7Yb8w1E
3KViUaV+wv6rYcLtMgq5Mt157tVtlzJEHNRQBKYACtuDj8S0CrCyMAacl4b8gL1M
oPeUqfawVfehOVfcEGWVg1h5jm0kvH2DmxvcKDUUUdWYwh7saKB25KOASll4wRI1
rqyVxxNUp9nhJs8Bjc8WSRStm8hSu69Bu470HdrilMe5rYUHsrAQ4G5Ye+E22ce6
msjAlV2uUi/SxBHK30Wfk6xTxeQwOk++P3ceB+KFLZq6Jc5Xb2CehCKZu04gIIHe
akPR7DtpN/IaovE3iOwBHJD3yErtfSGLDN8trWMrZ1/Y9se1tJoG0kU8NWWVB42L
TM3yPT5mpqY3j+125G3jtNUV5CFs3MKzrBR0hm6wLOie4Xq7f/pd29YWtzUFeixe
EkFrf8wnlewQXSKnazR0FabQn7xVOhkHV6o2kyZZMRKNs5aj3dH0NRZHck2R/FuD
owwucJaLLpW7YL3ZjsHdquhGH4P2ZS1bp/GWLkga1VLK6fXQVAwl7tVISIpQupOi
QB1d/MOV3vinAK2ZD6nYEylrrdMsK8m1jVI3yfcdh0hgj3rEQjlUCFI9awlHdQlh
hnf9/5MTMn5pnddmNwhiNCXJOqcKh+CtD/IFG/Gl0RUUw4/uHdGVEcEHk/CBUXIQ
WpR+IdnwTgQsQcCzSPcmrYWVkXBHCHLRuV9/24ukxYTtjhUu1CsG5UVieTJ6oqZU
vsRZOC8wckbdijuQSiQ6IFKub8OGEvdkjnR3KGRlaPmQJr2LCys0CWzTGXYAV6OK
EooJ0TjVCo4PmYst+Vx2Xc0HKkYTRtx4Z5ynx1fwreU4+NM0K241An7oTd6QDeq7
7jnet47i3qqgsIX48JVqSElNYt0JAQkm56gKyt9x93He5bt+yqcIUsDYlt3iDG38
4IwmliWyt9gDmxEIH6Q5gObvILvKE/Q2EQxCa66U2en1FGupUdvt8OWOwuCBnEv8
dln/4i/tERZr8cgI+qcOSVGAOA4226zRekS8TRc+SU74prJfn98bDObJATrgv49P
kTk9mC9hhY0tk95I0qNe3Y0hXkGewoT3GdZHW38h04J+81wbsTRrqmscYaKa0mcs
thgQ6XVbaCQWcmltFDmwxMq3xYej1q3K+x9NozEbuFtITBdhVy/x/Z75k2wZQbaW
aMZbphckJc02B3l5qJKzF7H2BLOxg5amlAkli0a2C7lX7eL3i7NItIUkrfgJqCxw
mcVnsy2BFtN6zKDuCp+DGHLzUgaYm24JTk5cHXGlyfsXvXLyf9VlI1MUJ73XbqwA
Z92tAtCmTAoYHnyOKQqMnLnet6fbOvei74XThL0MhBUD1OJryF3PZrhrTDDlSB3G
kdMDKL5OSc8edwCR5hDLQG/Ny4A2+gCtqDAAELg87ZPWQZEBJYkt2OA+zSdb/oOU
F3C1H45Eh3crx2j/RNW8ASnYPoBCz46N+jTDNbDdqXMk/Km6TsLRQQqipZc8rcZG
7ci41xSN7bVjEif1X5dnL1GanUGIknJDAkX8vgpkSUAJuy8y8P0nYXQQCUmFgpqK
JiSt3SJY/XMzCxrtdAB9FeeOz6j8A5nBoQpmGILExE+FSOJ7H95NbpYDw+TwiVgz
8ZUDEUF27adQO9Sn5DlgeO/xOODnwiSuQUFUUBamDq87xiQkOt2DLPg5+OVlNRWp
NVyKg4sT8NFg9mcTvIRcV+6r+/GEA7atf2hbsfX+imc0zJUb5mR3gUN1oHPnJlyc
ELVw0M6eIQ1h6lWYUhSOoZd1b74SEqkJP9k/BfDHrd2biavGvihMRtFQ5IcTImJr
xSsQIXLucrguEg+EvjuTn0d+PK2iKkMa2x3WH1qLwHV0dHAgG1jji1Wn340/EDld
oR3CpgvOrzie9uqYCvfYK/sEKNpqerShVgH3fo4mkzb4ypcyDh6E6MIU8ZV6rIUN
a+BizPnjUHseD5VPfTisIWGQ4aaIxylUAVzMReRc0Y5bNfff/dbvwX+TucbTzDR6
Se7Xzfe86OpGaKwGWMkqXZqoyzhr1vP66v82AbzcbGix3HUQchuLMcOug2eZWIt1
POnjfsjYtXUXAo5pjVfyCWdPLcMOjV+2aLdhyvcysrgk71IAIWhaSdnxLXe5SNyg
1SeXOMC8WCSK14TEKrBkrtbqN4Vj6pNhAFcK3uNbtPU1/fFqyKUkSP/LziZ/nYYL
pCSmA3IllFnm1k25UGWPwXKniiroJSuXaexSL4bzCesLXeKbxMtFg4Hb1HS41b6+
okXykpC/y+C+QoSb0CETPA3B49wbDKqiiZAm+VN6ex6FZlyRvfO/n7AYQTlwpLES
jHYcUf0mAjp0z4DUcfoL1IJW9kmvKE+9fVmUtYbnRGjCxNcbNiCLwNzGcj6kdSIJ
w99OmrTX6IvwSrOtHSH/34k39KQSCnJKkyEpMSDUscZU3MTtz0xT0Th4Bo5zuF6A
ulXPBBGduJXGvF+7vsWqHrMBiE53Dcc0KtLxMMKz/Dsh6X0hju6us2E3+i5J5Xne
jOuDhBz10/FDvPD2T54jxldSaLV1ca9L8jdQz5+neMg7NHzcL99y14PaXfBH70Oc
DY5gVCWnxk6dWyLv2j6haR07RHi4BZvd9iocTAMNZYIT3aCWlI70+zLOzyaIzwbH
xD672NF2ycRPvusK8N2ysmOXppSzN9OGoVNU97JgLkp4fB3ejvLpPUfd5x3YFaiJ
98Yc7xsy/42bd0wn6PoEJpKSo+X3g4RbbkMTAiKTHrZsKJVy8+oiiMRS/1rGofN8
Q/LC9r/zWHZ7Ut5PrOifM/mAiQsoY1OcLAOCemajFJ6+O9Kwf9aOO9NnJsuTnsl4
Ei9NoyNFfDndTon768NN0iEl8B9Z2ikZK8AIg2qW0s79+olp1sF+T/iW7ZjDJ7KT
dNudC8KNeMPgXpC5ny9ZIHz2u/5ZnRBiNORD15KesPpExd7bMLgE08vhRpxNoQ00
EjUdjWpJB9I8xvoTU84iZyRUPJDvOZphrkp12DkSWEVK10O+bOX7usTFXJJq8l8F
cRTtt/5rlnn3iMFtnAaxC16EnQl7EhDILXN+JBWbxPkPwgEg3Mgvxg6FgD8s0Fcn
DHymlPQuKEJfgUxfNRP+SJg32+f8prm/h4E9XDKDNrcx+CdKvOJoeVE6auOA8Ni+
llTH8Ss85TW5V2lVexIh7l7Pg29+0MwMu5epLDHzoOypWKwKlZ+9tr764d5wHcf0
4ERm8rUkzy8PEQ/SUrA0IBY5bLoDIwKFJZwob7J9d4Fs2V4sIr2QpOiVBTSe+Ohu
e5tKntYxIOIAa4Nnymf+o5zC5SEknYErzIL4fdw82t8kACeIHVMpvtTOKzTR2xh6
6iHsXQRDyVAox4KIJQUZDpwQ4AbDasXkBNwgo0WU0nKRc3fy8jMWUFdiiFpTe31i
twsTQWXhpIz3WoR29Cp+8L3a1qkIaGh3triQ7K650HJUsDqTKe9NLbDp3aKruUEv
NRpNP3I54BI3OlXW1UgeOQ8aYt3iObGCSuwPkdsCvEO+UqASHzX3JjfW0B6ywphe
oSxDaeC0g9mFIvVJHUiB+pm2vLuazCngsfh71FPA+B6ZkpCeq2JTI0UNi7kUy3D+
gjjavpoYQmLOnkvefd1eFbnK01gb/C3jEa70xsKY9SjI05YDn6sbjrkgtByg+YkL
zCGW/rjHSdcHeVHXuyEpFImu5Kz+R3GwlBAvsYPYcJmVSDgs/zz8XAb3n35b0yxQ
HEl7BKVKRKsjOk6z07g2pTxqN/aEollF3eaLxNkxOkJ0GL30tk+VD3HQzafHZIqr
uaFtfl34o2iG5jMjZJlrDhvcsMIgUvjyZEzdOzTJq3c3na9gJ9ETEeXTxPpeCBZL
lObYFAU+4k1ZZxXWEY6wm7vd+SmOzsc9daaSFis4NRqXUWDiEMgFlE+xcUcUAurW
dUjrXqfXBcDQuDrS4h1wzw1Twf+c9khLaK5tre3+sASPrVSIzrhDvcc76B4IIfQ8
E0SNNqAPWNDR9BLL5DkXvjgHK4+ccOHXRxZOFGVurZbLEp4lEbP1PZXPf6rEM1rl
7j/KDptM6BBjSScpkh0HhsMxr98R+mgZjlGUtF6ltvgekt5i+w7ksM9iKXQSSFIA
LkLeiCkviZnWuvn6iOFxtlszgh+Q/5x6XyhouqkyikwPOWX37zPwbe56h+AyjQEK
D7Nk/drA7VnfBpbK0EWI1LgOSwLWjkH6m7h3FzeNXliuv3VTZGabui7T+SHFrpk8
DfNxBoehXCU5xjhiJx7egQ/1eSkI37rccqpTBruggDcRs95pZEZ1Abqj/aMmMOnL
Kt/HcPZ9fyHe9zWx6sJDdeNSrn8chOJw/8jY+nQ4Iw7niJtaEglBsS5S0xkffxb3
7tSJsOEj3+nloiyG5gmxP1LC2XKraf9t63qZE3ZVrAn3PvvI1y85REdr28IwXZja
Pa7VWqBcgASgQTdUTXdIgj3JPwcx3NOh7ASHPgvk0zceQMcJxD542MJloe1L167R
A/kBv1q2HhpVJe0qjXb8ZkMWAODdQf+/mcuTJ8aVInnwlsytBLmQmHmYx2zR7l32
24omooYxK2/D1TQp+vU1jjfL9kuc58upU5oltouM99sd17FXa8JOd5nRo8RVssZI
Y5IOMndDWZ52v6OcLn17LYntLLx/De3ALU14nUcLZGUMe+FY6DDegUUF53gLTddD
SwRFH8BDJg/xZQmYis873iecZFVAmboVMPmB3wBHADt/p+opxTBZyG2d7fZYuWbb
R1JinR6dlrDdrC2IgP4AlKvUlBlCW6W2O1Ne5F3IaU6z6qzvNmz3udY30NfuQo8X
Km08YWDsqseXnSdjkXkHazrg+jKnAH7DdDOi3br+mzxkCzkzha/YtFKRP++xzg4H
iUKuZojzwqv8YdH4aA90dhLAY7e6LFami6yr7ZaUSReuVFZEAL5qnuXr6HILQDx0
Hq0RJuA6zE9NUFjVS67DxX/XnL/0wXPBuWo1yGpdSANS1b5xZWhGIzdNmPvtRWn3
jQij35xC0yMV9JFQBaoGTmbIBXYxzacsAbEY/Q47kNQF7Wer/QRAYVat/9bDEKdV
0nrq3mpL2ER1SKOJfHKAP6lcParFhw5xGhmh6CGOuN7fNCS0ASURhiTiwt2yQgsc
FubXGZFcfnqMSxoTu5N5zjnH+Jij4owB2i5KccJzo13EuPbt64WAoFHCP4Fip4mJ
a7isBOv0LHKzjbxqC+9hn44W2GLncZdP1J64NyHoYgLN5vkbcCVTXAFEnhypqjnS
fXVpeKQouHBpyH40bxQL/a3dw0dPXW3QAlbrrf8oINDUjfC5e3/3EQ88UDw3dHx8
dc3FgAjlGWbDnzJh2Fjn5mNg11HM6SXlg8M32CNfQXrvvW+fYmEIJ4WZCVlHBjjE
FSC7WV9eBf2JMeju8vrGc35BHKP8+qLdWf8zQj0YVCV++ZsD0nEJ+i2uAfqEdJNG
/gE9Q9OBJgeSuqFSHzAqWDZUqSU6y3GtALh14jQvS+Q8n3TN4N3eXxc39QIJZNUt
ISzQSYB7/XBJWoSf+6VYZ769GdVU1NGOsKRUnoVdFNDA4QfL51Ns12iIERgY8nwg
O7WgdhXkfJQKDEKTRlR494vIcCrfzBPQl3ryIohafmHipE4wMH8MuudBxArO+Zmx
aAPCFZu0zKlelwbA68xhXs0i0maDlNewntUQzOjkl92As5CIUr9yJQ+fnnjQhOcs
FtC3dyBY5sY0cK0X9EHGa+8oXIhnHqPFF4Xt7aTgGEG0sPDUwIxsOO513tBwiCqb
eb3jRSMM3WhA3Aa2EoxwRRxMXT4E6PzXUIXOFwfGDuyOWlBcSfZg+BLpXebs8et8
xolyLGv0ndt2OLThLmbfMRKTbjB1ubrbUu3LeMg+t2C5ORX8UmyDhpZ12/vb4Qyt
ZMIZCOAnAHVj8cIqkBmeIFC4IaRk0npMqbN1u5rqofH96NCAnSazgNK3NiB8lR28
YkPLv5ufY1sChEMLoD9dPdqCAFFHHEVEtiYGFwq6B71wPAAZzP9xnJ+dmxJXtWgd
uEfSBju7awF0upwPxcJW/PnjqW5BKeABGSS9Ah0tX/OzIcmpx75QFM4EBgFk7bBF
4y4oBUSvCoAAQAn39YwJmvfjCjYuaIi7HaKUJ2cpcQaJyTeR7TOR+mySv8q26rsA
x17XSrzIfbBULkichfFAQ0o74pw4m8NoI3TCbAdWUok0Uijo0Y+w4vNOixJbA+a1
s/x3JEiBbgVRqQHlrsYr+42v/W0rOeBA3QNCiUNfv8ncPDLxzb+Z+ClYvxCCeeou
/6N3wLrk5d/7e5wXadLJUhD43r7qSXkaSAelDfyN1aItZPk0JICn2Tqn/jk+ANO7
hsypB1foFKzu79ZvT+kTCeMDOTN92bWz644DQ0UdvjP8Y6e2FGp3wiw15r+iHCP0
zjPHwrJF8yCxuV6ed+2gjq0qfHZW3lhmzua+MlJ8nR87F+cD1FUE+r004bVOnW6v
wMGu8wL5xnzXLC0Jw1gDEiTP52l/RqoiTiopYbZBYmp42Im/T8G4KuOiyPKcEbYr
sX0UXTN0tXh1vwo3duZ8TGwE+N+807bRxx4jq6Pdajfmnq8mpDFG0EVkTu435I0t
ZurE9/+f0WSXI+r8Do7IyQZ4o4JalYTl7eBA7rz2+OX2gpIKuMDDdEn55CRp76HC
9aFnj7XG/X5CN82OFp8ftX4657KPN77cSx+F9lUvmQWigIjncXBOwoRyoPOaO8oU
aAOZqZP1HnJtn0e8NdfA3jjFGrRMqw7S0llniT66c8SbRv34NKn6pVtjSkzKQR8f
DuNOonvbxkM4gsD1QKCWbcwmxy4SkBlr9XIsHb4iXTCVSiFqK6+lGAH319Wyamvg
DhP+3l6hKoiqHjvRYpNuX/szecuqB/kcoYXAA6en3dAz4wIoWzdfB5aRVH1Kz/Rx
09vdzd8aKypFxM3pg5NyJnTiUdkH9wQausLUndZMMD+y5SYQytqAWwrOKVi8U+di
acvXEOSlrQd3qEYz/i7wx+sextHMk2TO+MVwV0U0sox6d6iWvms9sMBgV0uu4HB/
DRtKtIjiAz1kWaMqKbkh1bst8HFdhkYWp0O9sYtlkQPkg/ao0Fbhd273VWx8IpOl
OzvTtZpqtMtzs4EYmsu7Rp4TbzGI6mrLzqPcIL/tFbJiE3l2xjWYtJhfDmKOWPN5
Jwiw8fS/dDPPu5i1gMoynYXipp3eG7mOdE0MS1TL9dkWJutM4g1xZIrPQ1k5vlug
15BLGaYf+hp8sevU5cP79VuNkKOxqVNs8HT9iSfC7Jpj/iIy/v2sXKzLtY+iKYfH
Grkl1JxNp7OwAbLgSaSWZ3FqQL8Se/BevTxWKtaTWhTlb4GgqPs84dZWJi1Jior+
DrNHyvoVdaB8XLcb8hOdvy7ixA7y9aIul7BUulLLHgytAnVhKQYwcPMSENHhc3Jy
O0dRW64ORf1XMfhFBKBF0naPlUd/wQRdCmhsLYD11XvEToRPqDf1t84wOG4IBNZA
k+qLc9oIG/BVhm1m8TvTHRBpq4A7PBUCMfnLu4NBJhM4hjRrm+w744EPyuJx/VzA
/E7tuyasUj9OGbCzY1NkHEf11gh39fHIKXlXpiEDITmW36rRqJeLbdQuhn4Dzowm
tuOXeapDK3KaRLVKr+CV5hqRwe3R8vxSE4D7agATxcKMm3c5m6H5X9owZhRG9OZ1
ApkDCTRy+cH3va5uE50zwLsr90128fjHPpim9QyCNadxE5Y6SaZLVVurp6j5aJub
9UlclZZ7+m9t+5Q8Ra7r7pYh/zU2UGBYC4R+/RfqPoiDE0cguMVBNMENxmbc8csz
vzID5PGTc2Y2SwyxOll21iNMDV3rxs7FJjbbTQ6JcAX0If9iAwJYvsBRHrfbMJlB
ioTLjEvZ8AFpoM3wZhxVLS4e645gGSsm1mb0lxQW0sV8e8dpOAR5K2vweKk79SBG
BaPaeu5dpQqVGd5N8uHyUp36+ZptEvY9J9GOS+eAzYMRxHdUGheuxqScWR6BpaLK
YfAmKH9NV2QSp/XvMtpPq5Txymdr54krC7U5QZYMwa7oS6bPO2NZ3Pt3CNPhr79W
Fm7BIW4HnCtim/pzP1KwQ5xOCTgtGzguqOs6nnia7H6iBDPaz7/v/wAwR+UNQydm
/bq+HfyYTXDzh4x2PlcOgNevtHt0GSlKMpwiNUD/6TeGxNVTkWEQbIWcQbfsrE8Z
oGl6XTXQ7OpA1gFHluLz6n5gW1XJytuDd5qjANjef0tFKTKHupUYEoWxk3OF/O07
AgtLTPcX6KeYDtwoYq7lc7/i4V+9twvvdGyij4QTk9aXw1suf8mo5Btz00af0LkL
eervAUbaDBftAK8bS16B1iJu7oxTpD3BrggEfmgiC9TP9lq8BPeJKv6kGJmMgMfP
p9MsMICHRMk/BghiYsdZBrMdBn+LX31uVwbCM0xAv+3/uboP7xfQY1HT4IhUYXZb
kzOE840WMb8SedImlKX7ussBo6SDWPLmOCROrL5G84lakewzh43XbiR5JWVzK/qv
rLl8D4Md3fWvuLQ6E+7m9015fNyyrLXIP2clFAEqQl8d/pm61WuI33twEx/DtWD/
NArAfOsAWl88yIvhyVeqcHonk0BG5JXBwSxry0Db7MiexBIwbT6bZD5yVMYbANxM
8dBJZcBMVLuvaVgeR4IlKu5g4oh/xkykB0ryP9boy+Mucs/3lcrMVWG3Ta2zeUbp
udoZY0D5+fXynCUI8/u6A/Z9Nwz18LvmqQncBYcRPF32QgDpHpPcVRnzW+CEbbTE
CgcGtLyctQ+q/XugCsRIYzRap+ndvMwXk/t4Oks0t910DCe/jJZH+dosqBmafkaD
Lp9kJvKYgmHNSqX4YGy/vOA9DyL5Cz5sR6kh6O4QGDjsvp8XPlkXAqRllQkJjf1d
bqamVjoaJF6yuiO4EDZeMZ17BgZfQ8FiekHoZJfwBaiG686YeSwKcbktIoIveAaJ
aOsxB+WnsjfoqpaufywvzEtWSqKg9o7/rMdnv2RUkt050UxxYfjeo1gpXClMNfhg
6XD2Ecu1QjoNsrdYefqnyuyqDziWsQFNSZh2BlQFpCX1YwFFrzquO5qrC/WpgX/r
RRdZkriMqgbw6mbDsW4ZE9klsaD7ywa3eJmQ379TCqmrwC6sQ4WVp3c3iaTc9QVZ
pEUTY8tqTd386UhAyoqk7LOLl4zo5MY35CQFvG8j7J3MdlRUEPnLX8ncuijGAONV
swLl0oZVYla2zgBWsq0h05+yUKjrlYih5koFfEBkSZRv3Q6iUk4WGmliYoqhxvpq
igotGWpGkLCzpmiqVV/HumpaPtciPHxwVu0kkvKgCGO5owz1NfBSRmAIqW7ouTw7
p8bMUkbOWttmgIiZFtrCJ3IYBSa7R2BVktHM4e404AyuZmkQBgQf2DJWmvjh0kyQ
K92HtvDVDHO5QBNLrKINr5iGyfZGRV33BjBgKEkr9FBuaufqbShvy1TNi9lSHkjg
DkK+grXCGzgyR7BFIY29XVHyffQQMsSczK+q9J/DU9JlmycwezYWOBH8NG61ZRjV
1U2M0BzncLdGjUInUoCqG1IIQonXUGVx6R+PtlH/EAZpGatA+Au7JYC5C1T6j7jG
ukd+JEtJR6T57OriR/DdgEgH0AnqhnyC8+utrRqKLFtXlVslQMDjt9ONW9U08ob5
KdvxfWe5RJ4tQ8ZIs7EQKnPuUviTuwIh3yVp1D/r1C/eviKRHi9pw8j1ONRZvhUy
qUP1SjoifCpyVt1eE/UPQY5NxwDR0/bwtY3yICZ56ug+R0XNMNrbcqvpGujex6zd
LShxgvN/6gmDju7TmWTe/8QAHSepphykyvGahjCBbTQwbMhLM3EkSu/Ezvrjj+ag
au7tPq06Tufk0PUnry0pNMgX0x0NJsbeiqYgeTPjjg+hSotOU5RI702ms7f/3eZf
SHiUxMDqcso0ukwDXcHDlhKBEDylaPApXjKwTDxqvqdBmVzs3zJ9wpjkcnWux9J2
/2NfQypdUgGFGRd+7j7X2W30YQrNhsR8AvYpIHEC/EwqKtOiiLIomRv21YMHSBON
ecb4Y133PGFSruAG3ga89okelFKb+R2AIPbISL2lkVHjMNCcyoOVRevZn1VDijVp
ppULAFPySdEtqR1qgBRTykIzU5aS1shKWg+q52ZdWU1eHVm1CrEhbCTwXPlcnnMn
9RTNRtCUzzHocCN3cotHQNBPgxinLItcZ53SfI9KUvqws3VfMs/UC1aUPxSsrZRU
51EW3Aepk0QLVuYluphy+gH39wU2C9tLlpyzRf562kfOtLb0jk3XycojFMH+EkiB
r2BBE7gOcTMa9CFTou177YBBLn3tBUuLnmWr0PO3QvRS1MQuoyfILjjkMO5c4xzz
rzMhxXYphsMeI+k17MWn+fVK9y69uRrgqb4mUbpkBCOBZzGDE6GGOFugAW48sPyl
clQ8s0qv7S9ezSN95PjvV7lHjHj11X9Kt4Sj7sbFWoClNgoTu/c+v06kr24aVfPL
lfThf44r+4belQWEzILyPSnyWy1ZmE8ielbM6pJylxxDJCyqwVSboCGzfg39Lm43
66QfUN4WAqlq3PbLqj4QGta01M8V4CYxJpPH6UjhaXjcYcqX6ZII9cwAyfkSPTTV
G3eYnnFvkfrxb+WUk/EOj0l5XTKcyC6ascy3p/vAX9+e3Ui3HYMRHwXDtLFN37bu
pZ/owlwtI+GRexrMbInhzGRhoYmkhCPG5d6k7W8kz6kJKAUIEdMUC2YS9ZLtsPHc
rMx+8Ze8U4AqmzjUehOoO07iyZ/B3nlsnuvVkpNCx27e4HzfRYbM46MZ9skMKxyE
7gspyafn/otLZ/0CKRpocFW2ICWrOG2/BW61JPZAjiGYgL0P8N5zuzb77Ompw6O7
PcZZJYWMYH9SqL7d25IrHl8Y1Z9Lv01fKvbnkcSHSOAiM4Cjv7PXW7yEoWMBt38u
O3AB6NPswKm9mFOt7reR2NeFfRkyw5H9fULVIXlggTjqdhtp/MUTRe/DSxLYdeQM
g9YB3dJFuoA1sQcWKlFdlJoDoX1SNoY5uxsu0DXEbyDeGkEZmgIJbGMg4JMecQ9z
LP16gaNbw052RSr+9G2KLyfhuivwCqc96plhafG5KhgBlOT8Fr38+Akmljrc97Qx
AqJJ6KhfG3mSg7hWvTac0DDpruApfe2zwsUA5/T1tY9UcgGLBXc4hqZINvnqK7vl
jNZEvI9NklDkcSMNZha1CIHVNKmYQKz3uKvXXyPtebDm558+3R6StOPlTizXw6lp
G7lVeQHxhnrwRsoLdYYDzoroAN6NMFXrUANnsEAf76tGO83Vjmfff0kzDCCbPohF
Z0ghmwCwe2XEfVV49GK5rdLrLYyBclY4TReDSa9PF3oGqznwbcEtheA9ozxGfa0o
fhqcyYA0yfMqALaGXfQGSyMuZ66/pEkR5VfH5a4KzET6ceAL0urWzfQl/F2VuN9K
6SX2iQf3hRUbN90hyCXe1Ixbj1Z8oJT6+VkKgyhKGa2lINpGekYOJG9JvFuNWFvU
mPN3/S3o01g0QCNomB+QyFtCPMmbuh84ckEdtxkfX6E0pU2fQlHrWwh0Sz/j2H+u
0aFRDraeZ3lKGFi8UNjta5EdqCf8E1VRtuK2WP1Bx19D39goQUB8TNoIWYkULxb/
VULamMTsGzucCK9vz9+ue9MjYO7CWL7LtVG/36esxHh5pobNHIeDrhS0Q1AyffTZ
sM+6daANnQL/IPX5KYcwbN45kBtUxr41qvshFgQ+qrgvYEFo4lreiILMN+ceaBGm
5u9FEvLiTtqBpuq+9/MAcKISI+MGRkyKh4nWtpgSfsfT32H+7oaMYR8MmG87R9vK
/4VX+vo+CyGKUQuQ2ssfyEVfPWmR5WaULsnwgxkDgMu0jCCGY1374sDcbsgXjwdo
u7GDyUXZ9AErw/NLoBnbN/BDW0ZPNPpuyvawOCgl/NxRZvC7qCq7BdcCK9ffyqF0
809FoZLhJW5pEAdgZvergtwMU3rXeVMqfmo3xZ8kvQ6EsyuGxVQriimLoicWypMY
u6jmTD43yT/Qm4/Iv70RexnLLUdCL5nle/EH21Nd+aNDV9f8EKhhowdmITLlD0lW
pAKGjUV3yhT2+ZJRuxHkyIODjlvFHegSXQbhWcISYjsEktnvrwrTktD+XRcHhBMV
m85ZwdAgpYxteMU+tkZjLRbfoM5oSlq7wHdvXzHihu/IQtgVLH2h4wHbXopN81ZG
dXNCBzsIdJyE3kcsDEHOaJdyaQeeRHU7e5bwBv7kJjmSTRG7efMLk70NUpkix/1y
5aV7kbnkpxD1QZDFzDheHSxIlXMOrul96GY9bFYNS/3ka3D+eG3lqpPcjeIBdl81
3cHsuL7hr+odUMX5RjCOked14mVdVApBcPUlJPmLatZeeivXAa/i01dCOgIIyaGW
KDuryp/XnYuuRAvL5ksFZhmekPqYGGjLRQA4JVk7UCX7uW0xkq77mPFaLB9atHqi
Wu7//4jvi8nmVrnLBuiLhfj7e7oUyWunvmOGglT7xUequ19aRxmkkEmhqegPC8dP
4KNaMxku3IFmZMnp7HphTWZiU00Gf86Jy1B8u8ymqBiyM5SAPOqTiTt0fXCHcA/e
nJDBOBG5Qp9V0KHn4DDLpMznR7nUfwweKvqTI5CAQJnaW4tvEdplmCE07xwq5Fmx
/Wh/d5T4uIUEFJBG4vOAwiiZ2/i3Hnbbwh2fT7el+HmpO2AXnR3Vuvup4FVAW4ng
H9sndUxrhO/2TRKUcRgpufW7UjT3cdNOsXDHvJ0att8HR6Mq1EI41yoOreuA/YNN
K3DOnfI1r3PZUo1WYkhMDzwP6hyyJIp496t1YNcKOno78loKcauFnKUrisWla7XH
dq9j333G3aqBk0Tx6TkYuZKgQKDAg26raZCaNWE535VIphwktG5UW4Tjh6NeYWQW
lWmlCQNdAyheURFi7paBRMLhFNsFSZEja9SqEu2GhSve6/7OMP+LSHB6MiLkStXE
XfJkw+bRIynzLYiqKiEof1FrRj1ghdLWo8DR4hdAv7Z+WS9ftmz9uaxhNrOxkjfp
4pIBEP28JVeMrSKr06Q8afYHBNb0DL7mRVC19uw8duM4rW76b7M7DsE8OqdCHZcq
9u9ibRnHgcHs0eMRzw7Pe/uChuw64YdVLTy1AoeXbFbuZ/xTGTDnB7Z3zhfjabBv
T95ON70cP17XCu4K0LAXxh+HaqmQH7VgcqN/kU5bMew4BSMEpMVVvWOVNdWyoib5
LInoJJvSmST3FtVh6T+95ZLkNQqpvI1AH4ENpbQQQq0dTEsyUn0++brwGlCqAa9k
XHHp6/w4QFvkcRMjASJLZTKWcIU+nOnb0lb6gn469hGT6BZDCe0u0NvvVIL8Y7ER
WjvElC09enKafQIhSSUmUDvkMqB6XywHm2Dnd7l5H5kTqrRjLp3CWuZNpbBDhL27
CuRwWFKpBCWbNgj70HNr2ULR/3FeHZuJp1BPfA3pivulGm3JURKRbgDhdEZq7Hxx
Wdj/rLTo4iBE7Vlh4CdzRbuMRbPL68wyn9JEj1OEhmU4R4SwrhLaAJdhEsO35U+h
khVHA8gwzSb+2WdNtj37lIWIs5Oa9dHPMsruff35ASpVT/xPyQWc01nB4FRnvt/b
SCyXXSOFnfA6Art0WB7LhfnPdeX4V+AVxV+J/worXjiu/EK4A+5zOkzTwASJnZDy
b/IwgDElwY0xAPGVmoFDogFGzNcRxWbbK7aL4RP5fXvVs3LgMJslAE2pg5Zeb+Fg
mg/XdnosWviTUV/1DBZSXDwKd8q0zNMaZrs/1c7EdL0pwTjWcqEghVQz4jOLXQLs
P8MUxKAB6rjBhwG1pTr6GbN6vxPpVNDtOQs4ZPkexJEtDmVlWQD0WKaEstKSd6eA
RbXgAXmyt0cQ5Ct2scX199UZiWnTZOeeLIX+IGRg08EgqqCvvmxO+7bMDIn1ip6p
x6WonQik2N01w4BTGUSFJJJdBdf8hL0reB9pKswrlPsNgn/UMOCMzhYqcM7XW2//
781utgmvXn4YOciMRRLjrCvQHZyguuXsEt7L0dP7TzeCHtVg4uM3H5ne5Yu71UcN
6W5CDIJFdMMMS5okkZNIZU1iyf18phQnJf4Xu71Ki6gQZkxdk5TAHbOBQ/tFA4GS
7v9EUZvwKOIPuPrzbZOvhT0C6D9saQnSzph/uyP9p+bsLZwL7J22obcsG6SbZv0J
qsuGf3f1jGARN5Ye+RHLb3x74f5+fXqUto7GMMhvUd1IkYfCtI3lNG9vtPV6vO4p
Np/HUT7BU1eAk+yywL5x7iaHJtQGRGrz48bjERUmTYNUVTgHoMqyvPLfRMvxBZj/
hhkygSCFiGSOwc6RooQU31MIQLeWF0Bwh/XOVXHoSbC+nsvmXkrnIM+12yEFjgVI
vI9u6ut5xoJ+gcymKYsYL3WguzFfmLabL9kkobgJR3sTK40oYZq1jlr2wbrtJCBR
dNWs2M9pht2fQAqa5n+OzGybWzZmnpNaqZzohYyrL+MWf+DKUF6LvLV9q0IuuNaB
N755CB3qpMR6i+bxsJnCx4t25SK20B8nJCgOUQw1b3CcC9X27Lze8PhxPrllHkbx
vkPtV/zUa2BiJQQBvU3NFEuHFr7BYkWBSmBivh2aatwJzCyngni+7gm8RMxQHaAi
ctxctBXkd2N2KKndZEHeUdAboRJeHMLD0k1lZjWH8Qw+bCU+tbpqMLyNlmwkBrDx
zLbKyvmHFJdT2m6OI1mhWO46/T5XS/1YiBscF0iMEuYoLrB7rABp7VBzmpWUpZQb
XALnSKhzmX5mI4Bcm4c2xiaZ88ivpsIskwSG23nutYWubF4fvZBplyFrkpo6sHBr
lRWUCJXkZJLiLWtmATQWe6RENwQ1I7dxVfH7q1pMgTWqC1KcSM7A9bbmgv7YZcZw
tZdpMjyMRwawpJMPgdrWPcVAkqDtLQg2HmH8N0XMPmiZ2gfklmtXvEqn9mDiADCq
an6FINak6lRYgzDy+gGDzBLuQpFjEtpRgKYczDV7J+4biZdBR/S2ZPCNUKXeyMfC
9G8t4/W5Nwli7dUZkcHm0/VFZL55wluM7mfRqTIhd1gx5+ewK122q5RqxBbF2ZOz
jkqsrttJcZZg+p73KH2EoPsWuU3JkNS0pVkO5271qndqll26iBN0eqc6XuENK8Kr
QQ7E974OTvIr4Y3p1AK/s1sZVHsOVTIXJ4kc1GAEmxovXeDqS74NBw6m+EsINQuS
WsLiGMUvTbV7LQYOWF3feuis4MMyubTpAuNVv8mkFhL3wHSyGzEOiEpqbRKINSQ0
hDctm7EyaE56pR1UfUqE7+YPwMgqX+WrX/Ybl7u5ImnzrbV8kudvZpZyVXxFpYNE
gfnG8dL4g7jZ6AB5dWO7ajRNmJMTJv49IrvSHNt7zt2vCKvdxQnVty6QqESyFowd
w68NUjn6Ri3n/WH43mMMj4kVd1eHLab7Qe33j9SA/y9V8j8UWC6TxF2JdCcYC9le
BmDZDB1gp00IOJ/KokkDIItsUjyBZbNSkmczaYesE1o+gBppa8F36YzcHl1IcDfZ
OLTho+fECqgL5zTsvUHkDlPPr7MIIzw9AKLmwHFIKcWOAxqBMNJ9RbeU51jtnU0E
yQvRaSBBvjdquo0TcTUqxSHIVTqnUpaZRYRrqkoU+RfSE6aVDVaqK0I3bZ5wmu9L
kNuqb6Vof/AwLyEewS1KLh7f3b63hAspVzip7vRQRT/gQ/pAiNGFMGpkHIkGErEG
g75QGefZKPhFZLFgomhfnoTnU4JH6gghsiiMpYJORTDiE2ZbYwlSNzNlC1ZRSYng
jUzZASRYR8YanI5vw8Fa4F8zjSBpjNKDJ58fJ1Bu/e/Aebe1nRpGG7jBOly+OIIK
/C97cD0Yqx2YEaqD3RwPNgA5LIEI9e6c0uvmKSIIhBLWD8zGZN8Hm0diq3S/4MgK
8VjhONEMeudqPc9S9CN0H4jA1WuiolThqnA+SCkq91+KoFR7BU/2IOZ30RIxQVq1
83LNPAsUcBeDSOONqlkTh3ft49TTi7RjU4SFy4BpglZhq74kvvwi2C+J5XbvaWEx
fPNKyAWaoOXLpTfbxqDx6uD5JhCL29REF34yoM+ANGloBFoX2OlaevUXb0HjFFjQ
pIdmEUC9kKRJSa/w1l0/EMr+MugNXyiZJ7V4dqT9Ti8eQVz17Lj+0FMy09NBfXRc
i5mDq6E46sS254iDLuDcF/Ej2uNiT2DqjEeKhUr7K0NB7U6W/sBnG1afFerSe4Gu
KfQ4v1ODuLFQexhFZo0j+SvKaSdqauDWa1qOWNMlDD8Xhb4J1xJm40nSPM+mS3A5
ZKu7OEKcUS+N9ORZ4UljP5MXgaynk1V0KIntDaLBv9KzTZNj0E+y7zA5UJeK4EQV
XF69msTplree+sXQDQwWfautCkuLmUeIx/yeR4SO9iXu24+nYXeIOk0iIrn6qGnS
3V3gXMIxUv0X0v3pZue0JIWslg/wt9gST6SVwk3pL1vTXlI76D8nhBl6cfLMQNBo
tyw1XGWOlZXao8i/KqQhrlWYGy9CwP/NXxvFGANoQcBW8JlaFl0SNZOkW3sCScZ/
SP+VuS/tV2zQbXKSewnzlRI8LoM4ioXoZ4S3vSdyeAqJ1SGUx318760rPcSyY/z8
VUxZIknhc52M22502N21AxvKDN97xjSHzXgikRQWmM0LpXGPlzmNdfRsfuSmfaDr
VNH9ui+p5bouLUHV8wZPatpJhWn5J3hXZI3psdl7Mx2uCYeg0vUlboHQURkxf7Pq
imlFvtT9SDZNWUq1XTFfjy5eK32SzywJimvo7GtO54SJLcWKhs9mGPPAXo6O9Bha
F7oNLIiFkkoncNMuTsMw7oZzZYqJ9JM21tFkG1+BAaGudIqpkcoL5aJIabOjYLSd
k89l1FBvs1Ue6LzEZ8UN1bCA91bRtypqceWupm277GnAGnskQMBHoaPEO3SpJ37f
S8OizJJ/kA6d0GTTzWeHtkV44Pu76wFo1SDYb7HPymLqEmQSe6dIOgE2fwrakkyJ
V1QkEm8fw5/sPKWgUD44j3hiUsej7NrJuBW2x87twPgLcRcvqCrxCBmEsRzXAL19
NxuTqHNogqVW09Cb/dE0E52/yiLJPKjHP8So2ItyZfOBlexPxS98v5IR1uiTuk+y
Jai91rm10lv5uVdGpU9+yYy40p99NOxcbIzsX1NwhURU4iN5s3oSURMnixEvEOo6
7nXMPeXN1id0QYQbbpOmHlBH7Ona/8hqEaIJOjSSsRL/ujCRQpCMtZ+93dsIjn1k
18bKOcGAvpTNs5RCUG9WzOFjw2G0SGfL52vIPvPSzZ5TiSSOD7gEAh+3eZpw19f8
QC5MX7HasEaZsa0NasE0cNUZ2exPDSVGEuXhVHuq90iN4ocQBmE/7xUSIhOR4T10
0pHtLUGHT/I44PCsOZI9IZh47Rh31xjMPoulZpRT4YqDzWy0cIeV6NWW9Zui4MOm
iBmx/4kp4In7EqMI+L2G5kZCLDB21z+4acQLXfQ5R5DF5/z2mcpt2/2zIVAWWenb
mcZqyW9yUIWAdXLt8Nvfl/9rY6ugtNIgCIP9SO8PLjVtx4lqtLNPiOrcO2r/9hRQ
2M3GW1X5UyrcI9k6PQrusDZGR6Hd9G34CKQpQyG8Gn8+nQ+uyHQFYbDm/GszErFL
Nvb+Rlu4WTC+2ySZiO6PdmvvBbnTfz7UXqQscNvAQ8AfsFHiTMTcjF11mhR+nARN
ouftfuQXyEvmT1CaFM6j85w9JCt8XfGiH/p5kdP3YS+iMSZs/fRFDacinLAZunvz
DgDpXUvSKbhLYgoVxGFCxjitt3Akxtt18PQFtrcfIIR9eo4UMdeteIWDfyqBkvlZ
7jr80fJlMkR8FUUF08K8TTxzpEB2VijfM/r5ZLcfULxTORLpGhYeYpnF61kzv/YP
aioFvsp2M5Yhr0cUWcD+6Jcr+XjJpID5VPO3l1c20zdHSWrgwHm8JNQE4XFlSCS0
yrqQIBSp9bh00+VxBsCrd+Cx9AKStOYE8OMMXeyNuCmWj4fAA0+nDDsa9pvevM2K
WR0alDm5gpbU7yOZasUgZ4bQ3fPs5AEwNRo8TnpWAC30j15JGriYmp2zJQsw3hgD
fmIHtQ6syeriK6c9143h6BcfV2Mg73ZNr23d3+gMFUyZnhv2pKNqfS09Wqsu0Fuk
cF895GeRTTlLGP8xx0jSaWJgquUyNn0ZPu/aKu8O2hKa1NqYdM29uDwiqUjguBZm
5HLS5dJ8UbpHI3/6w+20GmCUPcjnGiviVyI0uxeGbIZ7MGh2wcq00wq7vkEy+pqQ
WFPu0V4GpSUthgZglrwtEezWaSBaIyPUT9X58nTFVhu+nlKRkDr7S3CVg/vDapSR
cyjSIjeVIaQnHNDv1ZPpKNYErPBIj8M5lb3FddzvzHpbsJnFKOV1jGXRHntXT43l
6uQRHZTmJoQKt/jPjhq1I1lP0VedPMBpagskDVNJafFykTv2+8Aq2dw7vmrOgvOF
94M5ncFq00jlGNy17v6LpRWovUYCBWZFA763eSu+37dgr/2bULfCweuB6fUIAB5L
b9du/6zF7v3J7GlvermsPPsEEAvD/ZzTTpGCDV3+aSFFHyP+BzFj8AUhkZ1M+Mi1
oSB+4L741nLWyq+Q6nG1BIv69swg76tg1xHoExGOGROkwcMv8JuyAqROkQIHbIVk
3ZMglytx5DEay0mnJQkQITQq6dWLrrRkuUgpxfmD/bZ2zCR99NwVfmK0zaVN2pfV
E6XOU5TLbmnSpU9u2RnWtcAuulOjNQ87J8jd7vu5JBYWeSp21Qo4eD2NvdpdXn1C
fPKS0/p9EHXdEFzten3n/zZFKpajjhnOaV6D/1l79iSsKG4RQBeYethUw70E2miT
P+MWcB1UsQsVVjA9gy1Q9DxQN9Mn/5bZ8+e+fuBAkjIUuVCJ0lGHi9Vmz8cf4g5q
cd47ltItpxjKSrr9oPf8oTAVbHOVv5lXHtJ0EWpp/ZulRZb1YhBiRGnygIpyoJdr
iqhLSm7yKG74iGzBGutp/CbKQop9QKwzQ6ymkoTBDhcTNeUi4tq9baS3L9+OoPrs
cICl6QOjgbe06vyn8qSya+dvBUrQvDyQHoQ8SmWB6/uKC77C2MtB7fNQXXaiCvBA
e/IptWrMO3JJJJRy4nxEf1Wavcy7+1ER/UEzwtNYqIYuJGUg2SXih5F8cvC1fmRw
jEdjB32RxeyAOdW+l+ckUAfThfGScEykWtN933RhaBMFMWo0A0yFvVGumYj7/eVd
kT4JxBKYN5rNAUcDPS5xRW4jSQhiNpAy4e4Sjyr0+WNdq9TOn8SpNPzUEp5vq+XU
erEeaVzESqg14irJRROBvCZsKkQ/Bx8gKDI46bghWGlLH6BAF2poxR55NNAWeWwN
g5EntfrMB8oBcpvzNRybj3jcGI/sL6AJJ+aMWwCclHN336+O/TW36SsM6xZjMx8Z
5RknN49ek5UJSnitKXjvRFkk32/mWh48OcYNPdxUQlfe8AxLpeiJTFjtYr2wCAyG
cBq4sKlfFud8ELdzJhK/R5SrkB+AprJe8MlROxoton9QwI4S9TKGquOrp8YtJEmD
ry9SeKv2BRNbjVa2Ceb8M/hSuXryXv3utZjGE9vWkEcI6Xz/b0qt9R/vVE31skCh
D4NLIGjcfHNm0/EkKiispidxkfbOZzH3+Ky4KzA8+hWLr3Xt58ov+CUdQ79Drp4v
bGm+XcTfG1yZDza2IPGpeY8MyJGU6hu0jc3PozHzk5z8hsqshgvIuShgTL5uSFSn
Akq4wP7JC42uUS48K+VsUUdZWwxPRW4RsjNmgeIh1dOonUWIydNkyDPETLQjpJge
wwyk7ve281DIogqLirJJKHgMTVFaeZ8QJXJALaf3ojvnlyjWZV5e6DKs7aynEqZK
/+rdkb1Ayju83JX3A1dPiRZHe5Q4l9PVhDF3VBzRbIedBlNdqDl/RXttZTXWemgw
H33heK8ox78XcXk9l8kE1A3R8LIHbfGUX0pIu35L1Wyzi4PsqDwbOWz124MTmJou
S/GnrFvPFacMkM2QGiR+ODjJu0Q6eiwEjAFBYoQHcX7BK06UEnVBd/SOTiK4kQ4H
EYdL0K0ifPWapZDofW1rJSESBXZ/23kD5hLt223j/wTfppJWYQKSjmLCJK+033Ax
4J1/liwpInpUX2Fs4evf8L+1gprPtRbMiJ1F8BRCzhHZYixV9I+RsNcwz8UxSzEF
twjeUTiGOIemPtaGZTFjycVCiAkBiVNCAnVK0hWkyaTI9OyMzXgSr7VZ11SeVVAW
QSh1aRK+HlHbDUm8HkT2tBl5GYlpdPSw4fd7BPQPOCTNEZeH360x+gx5Ju+8wGt8
r52ASa74/xiMO0/UWBxiQQJZyVoHSfprtstzykWhNFDn5D+D4kgZIw+3BRCiRW2N
x23I7peJV+FXf8FVAT/5JlImdCh765hWgrumh+KiYO5GUEc56mA1UeCdA6etHvJQ
r16YbsHWlHJwV/N3v9E3cLrGrUMQKwREuah/tHj/Fwv6zSWH//KYM7HMwhQrwozI
cKLlDZpNxloQxjLOf46Zj00wYYzjE9dMJFlS9jVEJ6zqTqx5E23JSDV2+D0ahUky
rmMLIDj4KDywdaLqIxDOoP4ONN5K8cyYUTmNS4v0/ray7Jppk21Fd0VJi4XyKSk8
hlDujsp9LyiPVPT7iwzgx0oJGzD+hJKz9B/f19aD4+9q2aHKwz+IllmLXF6c4Ena
ktuK/HYhIMHgd9VJVj46Wc3pOWIAM6aIPrpdMeCXx/C8trhXNAQmPWuzYnYFjOA3
rqSDPKtqFJSMgiCy7cK2sIWLFo0C/2Bc/OcpAkRb2lb0iyL3NwyMF8ANlG6OszAE
/x8WwoF4u4xiac43O/smA+jTFU6L7/8a2lpz0MAXgC+C4RqAgrQxFCRJIIHvVSqS
5VBtikCAG5e5pRoSzMZX5qjj3Jaf7nfElwzL8IZDNVRtwrd12NKc71AbfQdbyy5k
CRmG1uZ3cI2po8msL0GZa2qYlNV97/+qOHJRF6zWsxmgqbAwenz1sIZV0ssBK5ne
avxobAqCGUX1C44rZQwjIj7+hHiG8IugP2gtCfqamhzuDUj+UbIwXYRLQArnY033
sZxyALlbi0uQ+z0z83adkSWPhRjMvMKDF+/1N4ggIkf0tRn+pJK59aCmjOc9k7Gu
gOus5pmsekUQR0Vq80KsXf5tpnHfXFvLJ5jVb4I8LBQGtPj1xqy9L7pqkADYKoLK
V10VShD+gCgF184tJGb96ypbQEBvw0vrXJBnxiepu+RvPD72E4rZUZxlJ9F4pUcF
7gyfl/8qsNwaDEuDsOWCHOvxZ43bZTi+ZXwZ7zXXsqoG5LeiU9DrE5AUMbZ5nhaF
opU8vufpWJKowoHhD61GoDsvZzAI1pn5RyoXkbLkYHMR1n6lWlnughp42M1ZCZbg
fOUVLXB74HRajRzfHbFY6udYm1oUAQJLY74RfcY+VqBzi0RrA1HqS1DrxrM84c/P
/waQgmG0hRZZUkrNXtR6sxYCtu9VnSmUWjSxM/tBdnlGZMZQVxWkhLwbjcGkOWcq
8+rkldnFB/Tdbb55lmLOWdra+Ru5y1SItD1CUuM2cN8VcRC0hiZFwSFzWGmtmP2v
Rt1NYURPPCDkN04kZ5vfy3UvddixBEqaKyz2Ed5vZA5wD/I8Ples8q6iC+njta8g
p834aDgREdPGemQ4dIiRTLDLn50eFZWl+nUOLFJ99+WOmJ7bIF09CP+5fPXtKTda
FNVKypz/3De01xRKyENAPWpF2IVBTOHogaSLoWBr1blICtmvXJmP6SDkLZq8SJKO
7RSvVHOLwg5X0AnFzXLCF8ElD5IGplOLZEDQGw52DwuPDahV/Hne1LwLHYy9N+IR
hvZzSZT6U3eIAIqlbeULvuFzlGDTRgr0FAuC7EPU+5BjieuThcV8TROvsav1Tip3
mh74W/z8P4YLhTGUJYvItdbBgoZ1B1VROfDGYtG1IL7AkWLyP/bVO/cCLIbLGfy9
roDv34fBI34aXZp2gzsWp6g/XqSIUw/m7DOGHtohIgHMWncpHQytRy8LKIUlrFVx
D8gAoekG61g0/XwpwSNQ207D8WUYReBp0F2g8n7Z81M1UwTpQoub5GpbVHJP15YU
owEFS8+hT+5IKfurNERoeKicSx6H+w6/1AxSu0aZomKgDHK85dcfXNkHU68hierA
hJ4vmT45ZexwWofeDnTNEfA1hDKIJTqlm6GrAT+0w3GsUPCKDiBiAAMW/lpWVoWB
1Ps2dZMic07MJ9Ji8hMmmvcfx7VtDfdiGZ1+iELKTOurvOWa511zQ47s5nRcmMzK
ahyshexeCDfOYW697Zlu6annOhdl1G3H/NLwBmyR6TQjhxieCSishPb9XzKqTtja
G/K/h0eXfgJ8YgLo5haZ5rjctEKiwB57WAxsWUVmuxKJbad6j12nvAsIoV1J2Q46
zop5U4Yz6Mk/gaczHQwFexeTScJj7RblAP2r4CTe4L35zacj9+2TlIqnJupZ9Jno
aHXRStuiBeF+yBX4ky46pNmgVe0HW2bJatSgd8VkF+jmiQCEAarZs7B6/e3dD7AS
28jD+MOGbYnj9kHalXrtpYMpLfFp89VGKCWHfkWo0So/iLSAB12nC0BLlU8T2Rx2
T9dUQxcKZPKRHP4aGSRwUIiWweYEbYy7U7XwCEj8swsjcDSnrV+nIeR/oz1JXGXL
FKS1Ce4CYmaP+eUBDLkfg9C9a1i8rHi2OFL6OI/qP5Wd/BGHJ4+4STUd9GwNyCJ0
8mPFUTBLGwkTKHw5/Hjc35YS7xIfixjwHauAKpIRJ4hzlh0c/+hMZneojhAqfDWA
9DSKeottf/ztOvMizdqTPwbvDv2TqW86LDP0ONwOJIDTR4DbRriV0zmRZaYMSgAv
Jot7qL6YRmLFfBL2YdYJ+djJAz/FkeMyAarlsc8O6/evMfjJadfx4dQk4rVQdIyV
pOP1U3ZgvDD0AtjlHpW8xFYqCoBh/abhEFen86ShgYOGmEf61j8RHoCw4fvaLhNo
U62YKIzSeC9PG7wjT9l0ixf75wEKcSZTb1g9OQ23c50IXePDQEmTFTZ0W/2C7+va
S+itzOyiNOwxADhsgmh5dgLIrr8YeAjglb5d1Fbrda+Q2B1OhjNRnoBQRfauGC0e
QKWI8uyOtAQ148kTpb3WC3okBGksJuk3WdCjmhpAqy9wnDXOGvBLtvB0GXuNGV2M
JRXYGFfwSo+ct5jwhaqmr8DOwjN/yxcQVnntVFutZwe+hgA/DJRK5nNzqECxc1So
slad55fDnXCirIHzCNXlcJTf0Cuk+POtmSbttXUfUYYPpLDf9lZ53z4MGI+TU2XM
i6sZQV6R25Howl3ZWBrL4tSiEvBkqgKvJjFFhyoon7VGf+gRHSnwmYphYHYR+27t
87CYKs1iuIgPKVjOUnuZzGitjQcocg/ZqoFhwI9xoSmTg0ZTKZB1MpszRhPMigut
lb6kZ9cf96jNs1DroS8RYfy/SBtL6UEF4pYWbJN/JcxRGQJhRXINGGDT+xDHoAOi
U06xrep4eq4ccvyTCcU6urQa3Jxgw601pi2z8FKDK8W+81NOixKi/5ikr/PPUDTt
vMMnMqoYxtnga7lzClLnm+mPjzxMGy62mcZ+ryqJdwORWQievBO8fi8y/dyDorOa
BIViu7fSBTwEEbFhijn8bN8u44HX0jR5D2H0WNcfNQsAzepJy4BhDbXVbpRMK6gX
Isb12Zcy5FVCCl/VSKgAKib/tORxG7NDUP7rOjGmsNDwiigjoRnKKzfKcNZ2OsYQ
4lHHZl+Il0hPg65KWegu0ewsHitDct5JwCK02CEXK9hsGKfNSCPiI/AeFO3mEBKn
qDuYboxdlHIEtZOECPTrFFLXea0cRKfGMS7PCSaZsB+l+G3c0Ie0legrh+4KcZr9
Mge2wGZGvSKC/t3ZneYQF3Q4NPhY1wsRvGjLFfCDeeNs8sz4XBPm+yqtFpbkmN1u
q/EtfkWb47u67GYZ4ZMUPVmgrELMLNvzkuWwi3c5j/W8EK7xo6H80VoinV1OUGJX
HvD3fCKcnTlLka6Y+27c9LhfYr1fM7BU6Bo23Ldq0O1LU0D9JDn1eP52xK90m9N/
S6rQ09WqZ0IbaoEE9rS23Vr2yrGqSts4oSTRnz2e30PFKzsl5Jn3uLoGWKWmGQzR
iEN+BI2PAWCcz585HdEKcXqgGZUOC7MTYmtQsFlxfDdXo8NVXemF4Un8sATRSbrw
xa+Nwrehv2IVwK4w/y3GaK/7kVe0hOYpMkdA1KbAarCO9yNftrIgQb1rFyQjKcpQ
C6auNPYZKuMab2+oAct9iVNGMndHT9QwyNJd/XjHVZ4kPMoF9gyJF9JaGPMJ9qou
1hFBSIOGn/TYcERpgvW2zdpb/l7fcJYGpY6E4zYXf9Vk+RHdkrOebKGK/li2lyAU
b9tXZ02NY1sEchEkfBbLFlZOOoQssfpvECrPPLTgLonBkyT0hnFdO3vTRRvo0m+B
fZYsVaXbJDHFapMgBtMTPJAPYP/orkmnmLEE0QD5KyrQU4DQWzkzKQp4nqfQymnO
GshvrdmxvASqXnOEb1p2Br31tYEyGHrYelfq4wQNS94mlYVlhir16trIiDX+uzhk
msJ3GeB2x3filNOqC6YEKnxKL5N68jFSlc0VjMqP3VCsEEOvDXZVANgOfaXxl0l4
SPuF6YZb4kmCt/G6W3Qf7qiu9cdoiKCr5hvHqWhoxnuUT/M6ADAHgLxl+YFkg/fp
dZolqzoXnTztQw+4rSgVhchkBKn/By4kCaW9AzBiS12iuUvUMySBxJ2dYnCIjlbK
ncLzmPzKoB3H8Syk2c52IEesbIL9tWaf/oBKvozmocajbmus1E9r6X2pO5TLUhI6
wUj4KiO2hvGpiv+iXDCDVUdpwTfqIK7xevj5Z8972w7r7eD8cFqY7CJc3in9shzF
6XFufaSnKXhMJNlvbNYxpbGK3de8BcvgeOgNKQF24rpcCvroKfYOl03mR0qrCthU
o/fp46eblOXQKotAUOyKP2LGAAKAX/Bgjc1ooi7AoZFDZyNevBJDhZEXgBgI+fSJ
0m/SUwDZqQ9agvHUwC6ffvTLcKvemEH/rHMrNztbr7wChIvL5z499XINubVxQZME
WRVYHUkf8v54dIhc9koDcDNnaUB3Z+sg901w6/ON5zghN+JT/ghOMWUEPTfgLnV+
RkmcW168xRjpBmCFTzap0DiWhE+V1hC1w/3JQBNzgSt3y9+VCat+SoPW998qjVSj
iJj9oSNmN6pGdAUfkePAqOUbkKhtflmV5knaRQr1lQCbG777WCt9sq4ikolYe2rv
E4WIESyWlogFSt275XUDd4Uo67LmLfu4KEpM2JibEyIisHa/f+jyiuvPeWaVqL9/
ZTds2VJNm2dWcGrGp1s5pU2OGSV+tu3V5nTwoHkCvJiZ7BDarMlMi3nfSeBaogqh
4p1M0wCWOnSU0GgXN09VTznJZVuCXUN7Ufc/nfu6F6eK1rPds2LuP+4LboZ/VuRV
kaqlbNOO58oUzQZxNhPN7VWQGXuAxxiGjvaWmZZfOo026QNSKaMbIpQWrWFEXNCI
98rdBVoHGzAYP+pTsPVI2tp2dbZSfeVCJvPiRM9yA8WQVozptyUfAPfg66OtSCws
YwThgLKczpuOtJrdMPsMFZ7ZxnXeWqp62EFfSJZrP9KZbtRYgEzLVcfKSytU5z+J
/bnEgmfiEYeIqLS9tNO4WrTvSzYcJk6vEyV3aGNC66EXLg4ahv+qrG12dtfo++yY
TBWHKuXVOtbjuOLu3A2JclDq+xvP9QYklIG2Y3Sd9aF4cqctQCet8NkkdPqkTNrx
33zHk7+Llr9HEhV1cqvl1EC2rFKFe/VkZnQGAyFbXzXW6fi5pD8n6CX/bjvRVbRw
0xvnM6TejbovllLHaZLGITHJ2DU7l/OGTriXeddrBxQ+NCTkINU0BqFks6eMhnXr
8+4OljfYVT0Hqe/eHrl6/yoaZvcm3WcVl947Pl9bjLTmN+vC9zqxgjpXWFPgJSaO
pyWIXavkb4M483uv4w/uHqrRlYkEedrC9B5gPPS38Mpibf87bvg87mJOJmsGXksY
M9bJgaqp6YRnrw0beelQM2NBUTFgW9DwlHw8Ry7ehnVfCab8tIBrjO0L+9hQeRXd
382Fk1n+5Pt/ucbq944Nke9SegJQPUIFahVTxTtvYz8oZfn+DbpiXE5kfsnYZUsr
rUwxehgB7iMrBEZVfZp+jmaB9YP6jWfc7If7gJTLSkhfZwlc8qb/HjsMUD/PXPxg
ZJG2/bgNHR2Kx6rCyQCNnVdl6WxPgwgLQ/m9lsRUGLQBDXZkD3ocd8Hht/qGxn0h
f5GuvxZE5826j/zeoDwRLClVU5sRQrneNjpo3dyZmat2raKy4StBCF81dGKmEfrM
bVBRn0ViYFZ/JSNgDfBr5hu6g05Ld9Hcnp499lNivKNgYapO3kWBWaJ1TPLBt1LK
0YDNjOIfC8XEpMEayvxVCRy94ELtMjPKLDW5id/ZHbMTcQ42Zrn7ryFR5C8PLvYw
wcbDc5THxrBxIJTzEVnwWQlx+w+dmynXJAjyOC/0jzrIlBdHiev9BJl1a0M7Sw46
9kx4yjRDrvYBiIv7Xf3VHc8x3N6YO/SLVv6C1Yro0N69AZzg8hiOo9zcVAww9VTY
k5ae2+gAX2F+CuroLprWhG+lEbtO6Sr0KlRXRv2Je+btjWr5XVc6CN0bRwEShPNq
wRJpHot8i0PxIZci2M0hGu9Hcfz4zK/oOWcqv+VyOgdFATfunKcbzY2vCA+Jse5e
x4OuYZ21VWgf5i/YBXWnrkh1u1VQuIYYlKX28vjNTSCAPBHGDOn4EkhoCQqfX/I7
oaRqg7Nxh94QuXzwJLOsS0VELGuGQUW00DEHk2LFo08R+jcxZ/3fbFgHYfJNFzij
dFIak+wOOaTJoEP05ioO8o1Hb4lo91vgyTFBwtf4OBc/K+mz8a0GOlJTtKT3h0RV
DLPSFQBGb9zNg/PFKKkI3w5d+adsvBl1N1MPkiT3uhae+kFa/s8JSbBVRKvvIS6x
fiTHuvzI0av45+l8gXBAPTFotSN99iG1BY4mib5bZjHQwmEC18ESf37BqmgeDt6Q
RCsrX4f+bGCEPPCeq27KcNnzIcBHbmZhsqsaplSKPBGRBEEDwLm8cDcxd3OnfzXo
7qgZVkbrKIB2XEWDxntVSFPxyQpyF8TEBJV5mrGFtp/9o76ORyp/ljgi/IDQr7go
GQP4Hla/0JYgcIB8Ms3wiPkrV7Bkqnv1MpLtrdj9wzmYbA0uh4zzvoYSYTxeJxHX
crJrXHfTz56n/R2oGrGWjBdfoA2NZGUEpnqOrjQoQoj9at+cE4CpFnhK0IQup+NH
smSU46bLu20yc/xGhuJ8GmQ3bX4QNKmBnUA+Ez6FMD84IAVdToVc6lSl4DWI/5Gw
ly4S5FhdoxNMcf1G8Doo/pLeV8rvcjyshH4e0ZbPHwimWXhkxOt+y3U4hhVdpqb7
mq6AeVheEGhiodos4hqsNrUwQy66dqE0+cz+yr6ErZ8tMRGltnXCP2FaDrcduMnV
J1mokgu9JQkSLTQKLEo44GgoEPGyv1Ve6CYS/JaHm1lCEiuMepEaT0dwx7OKCJ1u
yVtA/rEiu5S+68PND2Tx/Iq9Ya9qBTCTMexlosvXk7kIPwOxkCjjBUb1ASAydXfs
MtiIFDk/XMJQBtdxAa+3CV7rO0anD/sTFtV8BtdBidriSDVMWton7zZE5xZcwTYA
OSBeg9c27Vjh/7rgf+DG/pqH1N+ddXBPH0mlZ8dvNI7olQvyfffXwRmpGKTqe+9g
KezSAaoNB5SiVdAC+YGtgYVwcqMXQv+74qlZ27AxIzLJqplLtfZbOX7122/eUZyB
hyKADXhKWnnUh+w2DVhEyG9V/uTAutF1fXU4ha4z7hAmlXiLaidrL9jJHBmoYH8T
M+K14ugV/Oj3AXSXR8mVyy+sMpqU+pEqNJSjH38eCuQwQxc0VcYYfZzwgieUIwRF
VyoY77OoWXA74RTYUkYChZM3gZGNNJ+ie0SA9GHcJ1os6IMiu8JdMbUJ5cZlaLx1
pYgfseBV8ZSUir1aDzNdoV2BEcZvCcc0vdbug1Xi9kKxiYJt793cx75Fd81k4Y0Y
bO2RBWj6dYBWLV0Xm7VN0HAPG1oVNgnFWnpF6MWqBW6Rad+Gn9sXZDbFNlMn1tcv
9PcIRhafnFLEEndZZBDGOXMV9wyAhlBcO1ALke1hYCNAT1WxmovK9/M5+HMqLvxx
t8A4VtRQsPLK0oqoI6YO84EVN8V5ajTm5sDpeXN/8Nw3kEjsPeawU7tSwnDBGki5
rofaJVyhmx9MXyLQSLGpLckHm8rPbuYY95/6s5JK9APL7vGUoE0AttvZa4ME6ppI
kDL3uEP0yId3pyqHXqagNJrovs1w1+oIXkgMSb85mD7koRWv4X6hVItKbvCsyESh
3bLyxC6cB8JLrRYJ7ivs36GVz48trhx/3zLjBpyig0qJt4LRJ6V+PpItrQi5ZhB7
UkHaYmnAvdc7jBphCzhJiUIQTcUwa6VDKsc5r96nF2bLZIR3w0a61HO9IK3UcNYa
mdjQSWsRMslotRwTRlfu+vFbbLEKRY7EsAovRGUPJVPNtOlMU8c0hU4yrrOk+tc9
V1R/0J5n5rCPnZ8wo4L8iwFzQy4ofMD09s/wAoVNmvUww07ID15n4kZdqbMnjy9d
foUVxNZgj0/weasTG5sBx1DzYMvMg8bm5urly+EFtnAKEDfiaOoyE2M2tR902Lpm
clkxT/0tqrCfdk3x2gXvD0nePSqD4RQcFPB4ueMwCfsDj8xLXBEy7KeXFQ+0juir
477LYEUpLDnTI6CLeHNnW3tRdQogTwXQXPPwRuRlkLFHV7vU+VzEGjLHgvo5JPxl
HlxQ9ZrL3t2pHQdwyguahRz3of/M6xw6cqlnwY6uzkiyMUPx7hLdJfBipDZ3Juqi
QZcNf5nvakqdrsbJZwJfMZnXtjH8IhbKIV6nZUDXD6Lgs6oGiRYqQrbDn/1AKl2T
L0TFnbFhfHdWreWphe9D8L25Y0aMRCJFlJjoKvBbS/4q64RA8t6o7fUbhGkP9/8+
0Q/x/3GzGdupry8+HQxfcXqhXPDPCo7wDOcKzkuS+9Z88q/UBivqG5XOj/Fazm/z
zgxgmoxN9CqYw8Ce9vwKKTfMocXEXPxHOsMmIVFRR8Me5ZBQ/+C8tH8lBSXCR9Bj
H6ocbfQcfIH0FBe1jatyc0RjtlGQ5aLRPo/0mXlkhHBUCDZMq6CfCJ9SKLM7WbXt
B/fVTCHl1Xn6xmb97XxQEOLVbvc1ZCjMHLoEi6VhZLB5OR/SQ3y45nn3V9Bqx15S
DSHrDoMk3A8sAzk5SaSybu+zuzUXrwcrAIjFWKrCaKvLXwQJ/86d06NgAoh8W5aE
SO5aC2tRnPvdS36l7kd5xYxycbzwEe6GZLefK736dhqlZ7UilG/avo8ozPbnlxif
LGHDtAGSGKeoq8Vo1DaMTBFy66w1lXU7UQs/ZLsyAgWUuRD+eDNXR87WB6+tK/O7
yL5UtUptHtMl9SgrfVbAfzL4X7/RDibsAr6AXPmadKO4rPUVy/+KOYPWGosZoIfS
u/F0o60NXAn4WTxspGC+lnK6Vrjr6vcTgkv7WPmyFflwcFdynC6oxFsANoRwfEkZ
P941/gKAd0zN9pjrRwahzeUiX//yxMr7JgUr/tdqWwK8PW+L+vgjq4+vT1IJcHgr
5SzoqE+nlvV5PIEWMCtiLp+ubjXcZPe7eeOdjJEgra/oqlB7DOvfVSNxrVBs7ny9
/7l9HCPIqKOGgs12jLbbRMuOEyA/THD/ejw1QNJfkmlbXgdZqFFIdAWjRkqRr5yu
thQIKy71FEvS+HMNl3s+86BaLsQnZPLaWVQ/10SNh/l5nTkQURmyuU56uYrE0FY8
YFtWc5h1+QJYRDlb0Ic4RgsIimu7XoK1IxHAYJKMWvdy8LHCv9sbISLMw0PqC7NJ
fFqKo1VUmeaamCXy1g2jBbATUYJXhzBVV+ShkCjoFpbiBNLE+uN1HSvBtpmIpbdR
kfBqnRoX2jGwp6sxh1ovHjM+X5Pk3P8FxiddVOk3jhDtctkjCIwS4P9nX59GneNr
YRAVStGogW1vnyZDo8lRcqDkSMUGZZIRaSKM2xagxadm2tB5rAND2xciaBIxJUbE
UYwHO3atSS9Mvvfe3f8D+d8wg2sJL+4NNFqLgm/GJOwJ89CX7gOa2yROR7gnrQ8X
DFW6xc3PLnTfBzIjewOAWfS3bVXjQRa0+5+DlLIkHxffP/kusHE7gcGjhZ8YfpU2
HHq3hq8eML+8r8rj+If0CW74ppoVwly435mWrzCRjxRnixPNRlephOnBnx7IKCEN
s+vaWyDgRZpTjeYEm9xawquds5p1zoFovcCJpKYnZe6ZVFbWuCJN/+daenzwgZUa
RC/ckH9x6yuOqdEauFf+UuwAGA2AHGDXE8oDXoHui8gX6EQWOdNozzDTBqffqvTW
6k2iSzAC/CNnUw5n6LAsIuxJT2HWxlvy6SAeNMWYKgQc/K9wgByHPzPZykS6ZypS
sfsYY3O30Br3DZ/RcVmp3ws8d5D27kEnt1LPaA3iOjGPKbNDzWEQIYFkRx50Mv9B
M79896dysQp24Kmrt3I8W7FY/sOkjyToOB8CqOJziQyZhPxjpEp5qBUrMnNtyFsY
UUOWYReOM56a67NNze1AgyYQUa4PBTmjaw2YSCqH44MQsrYFEIH3yGqywK+jYX0q
Q0eRGHe2oMtD3GDTPIYBK9DVlIO83/YlxLGivjCOOjVVmKsBYuZvBcf/HA6ZEbhy
T8teAe7HJil7BKg87F6XDY41jwapH/c2aGobDRAdRcQ0A4ST0puKmLGHj+txaxrH
uAdJlrMFb1hvJj8NDkmo5Grd3IwDI2+BleZ7XUrpIzQ7dBMWVQ8fH4zLAhMed0hl
rFbj06PgTezWY/VdHemRgOJYdAERY7k6znSy5D1I3SxX3ncYagki7Rt7mrXEtUar
UZT7NaSb43VePTLItG3elcBH5pxND3GnvTz5xneI41x0i9Qd2r/Ru5L1g85ELFHk
2vyRYqYPIUIUXfqoQgEdkaSvDq4zZwp2/tveoJekf3Y0D7iye3KL0KHFeSnvr0WB
1eEoCc/1XFH1vfi0kffviK5SOyLBy/he9p8KGpVST+yqYd9/s7HzX2RbJSfz4QXh
8Po9WgQ+V3Vv9hEGZw529fBXEkGYBWHRkK0lA8pxLGNd1dqKMZwGitXPRC7416RQ
98Vdjh55ss0w+m0Hew8W8iND8d+53j+zIzsZ+hklyFhIZkBT1v6Mt7Fe1W0pjx9A
rUMit7T+LDI9f649dC11/L+CumbqxfWcW/ITrcU5X/o6skmdTgqmV3asHt/ZpS1v
0/nWntzeDYSWqoD2qZa/aO6Rl9wRlPlq6xXXsTnzYodBqHMaKIEF6Z2fclHEvKUc
ZWWZCtjJY/xwQvuvjfTJqtHS3TLKnFum1mzDm7rxBH4BJRGOUUk6VP0ybRfbZUTf
cJE/88VMsURXgVOI3fnzySjo7miSg9H8Qmq7n/xczEULH/JOm3acHguJ91a7SZHD
3QHothDDqDnXHITwfZT5tKgWTpbYuBp7jIuUwpKAR5FOWZHFJa9ty76PG8Sats5D
VVPg1Wt7Rp+BdcHfDsZMHnZlsAwRQyGCvzMFpX73fNLHT+CoimWs3lU2YL2d2g91
6K2RyNYXz0FOZN54zSffcGhEw7n9JR7gEf3N6Bl/E8TKIW7V5RcjSJhwk+xjJxkt
qn05LoWwPja8vaLBeB3tAiMS7Rxf5HfholavjBcF5aZOrInrWLRNCet1j0pQmM8d
BdZzZUECHRMxqDj6GB195xodLXNMM4fkvJO9blrfCZP5TTvnNw69HfAiAwhvOppq
qaSqm5uRkSeAX+tjTLRLn8LQjuGer6Ij2/sn6uDecDWvZU1opZRGwvtkNnt4oxF/
Bkbcgh0K0HP99MOltOp9UfeW0dukdkrTdGb6w/tJdJflk1ivTO6aLvvWLX9b4hQy
Qc5BPNswpO900W/BNaOafi7trfVoZwd12jfuEj8TFDEy5nl+m0QM1KV+OdYueUzd
bmN+Jq/2yj0sjCHrp5FmQcza7NjSBaPZGumdCFrQqpelx6SGbbTjcc3WezS00+11
Oe0s8ZuiT0UDpAcX6roa7Kh6nbeCFTgLNlWuw7sjiSfyTq5z9cwJ5hhYD8aomeUX
6/bpeV/n+TI5Or/y+7jyHUmNhCE8MVMMkQLzNvExahKyTTaDSKUT2EmLJom9M8sE
55R4mGlrbNxCIEb4rfo0slpKmPUyYBHFXIrfcssrSWaAJKq+3QGRCqyQZAkRU1jk
4HBGi2SmHijzg+jyT4HZTsCRqWhLGJM0L9uuJdGBwqHnqgfSa+Ei/8V2wJdlgkDp
6jEv3e2hPM5az7oGLQ+Gd/j9y8XgmDp/3oo1/mpgA7GXOfJ9rg/PKck+d7HAs5Xu
1ZXUEnasApO3ZJOvXFESs45PZ9v+jC9ZsfocV3JccwRxcO0VE3WefduNbGL3ssF1
GWRroBSSFbljf/1fU6YxOOBbLZZmXVUBRGWGFdjPbIyn6Slo7ZyAvr7s/Ujxm9xM
JYqctCjFBeuGmqVMBK7Gs+EAOFGgxnAzSsYRGPNxpTCr4dGp7Is85GOUyacda9Fc
NvV8FiEzL4nu1jZXgZke1rt5Bf9+kMUpw7QqE85pCBKNcjahLXSWFBGO9hDKJJxr
Eaqb08gukCvjM564iYnolwZpCpnYUAN+5L17Fpt82aCiol2bfMOYZWFw4jtKyTIY
QtK6Yv/oCnjbrfdDApCGzjD+fvIzI5D8b3w9XskoPKCUlkR9FhS0vmTCIy+RF3bM
22qVsECttKN57b9ydZj8EGhlTroXbGN1+7MejRdVQt7/KylxOKpfBoWmxKoYxBst
GGnaMXis2YWQWGXx+5x9ETitRxvIeVgdqzLPk47I3wmiulo3nL8h2XAy5k7a6Y1w
Y4dm2dVdGrT1KZRVhyArmpVavbLAdGgpAtxc+xIRB8E/q8nD+rmu1kNLO8lHOQqP
Iso9DgsfojIDSTHXZUdYMuwG7Bcos14pEsUU3VYB6JcycGsQVIVrT8j7ZcIqKC1s
6oA7iU5VJo3ogQjRcL5ye0Jc1y2ZOG4UJmF0TwTufSv3ZgCwwBJooe1orwlamJT9
SrVMM1comaYfGxVFvLt0P3t23D0Ob/mlpDucCKldL5xpqtc+tq54wxDouPuL05i6
mvLg+/C7iy7MjjZoGvZDpDwBd7SCrfR+5PpEmicl0O8y487IDgTr0nfLyeGSHEdM
JcOtW73Ytk8t7jIKx6CYQ1uCKSPactNEO/btUbLhRg2YPiFxwcWqQq4cepyJckAm
6mzfMHqyCqm5pk8jO5NeHdirA1V0JpSXPGs0utMVBk1XutAvm7bAIYikgdSLpELv
T2HASI+2zLRhWSDaqBpCmxTX/qHv4+/pE5UVr7s2M21BhELQwi6YRXQUCHMbh6CM
dxqOyRcasK9xrXwA6TXTy4gz3GA2UAOAPLo/IojP1aQ18zGzHOUKbgpBWGCvjazW
DNB9QrvnzDPFHsqKpMnAbuzdairnAmfrpkKqoQUlpUxOYqVEjiITqbzFEFkwbLiy
38ut+p0w559zsy/tjsDwET9WvIQTz09b7uAa5xCAI1v/pAp3x8iFLXHmAMBbk7nd
0p6YsDTR5H2gn0P7VgzNE1R37lyO/0cECDunwp9pjHAYgKdQANhBjGGKsyKRtjlY
/5Qbn1h/TjldPmnahfXsz10pt+wUasuURLjS+QbOE61sMwTXykyaXnJ9c1jqjg/R
uTTu/PXZ5aaAeHD5AWXnHRfeLnfaBExBLSabI1JkvgZVBTI9qgmFonwcis3SM2hS
m5DQgEwQmqMQhsdN4X6xW07MSAOuNzh5lTqlaixxaKlDW7hZQgIBEORwlZtvImws
xQDNK3io1/P9Ua2AsXRZA85Tycs8S/LRnXrvVTGSfRO6z+yIxiTEdpKX3wSSpH03
yAFk6jmShVEHLPLN5oj8FWUthLe7jK7CTZXWWHVh2WWW0G8igo95Bh8T+0t/x5ed
HKeWXMX14ALSRZGSgo0OyxFyNGzdl38BFnFFf1qgJbJXBb1qzcBx46i04aE8wnxn
bSfL9tGP5BWybFLo9QHEO+AdD1J6GxmsC1sQrjyjNF7LiMmmuXk3Ipv7v+67PDct
kBQ2af1m/S4DcF1oKAUD4oveICZSdhXzK/tCG6DCfDZo2MLplySmj15d4AWNbjAI
7tdZ1VzRKC1hw51sPddxMlv9/pA83+422kRRcgwlROnGATaEWhX2Mpp5OIFkLYNA
ebxphstgbmS5MvsS2Rqj5FammHpS2/o6bHQ9dhQsC7fLs42YPSMIQj/vTCJY72lm
GmPgt6xn+3/MgwU5QsKB3bn4oaw2quCTXoy/CrqaLQweYwrYQjJPU1eE00UfSsX3
dgmLaszj6f7RVnh2e2F6hvVD2ykCbH/9sTwjOrkvGm9+6weoTZpKzoxlnZUZGTKf
w6iZZqW8QyG/VvGDNaky3X3biNvqcVSgJYG3xsGfR7cPyqU3iSF8ODaF97//IEMr
Dsx9KrpiVl24Sj9PQCb5j+rkMps4gS5dbhDxEWz1RINeJ/Z7WY9PxsjRRpUWoAbo
FIFlUeOuNwHewCbrEt0PVqbCMv4Ljy+oy/SA0qjyH1JE9byWiYp0vGcF6OcdB7pg
sisG0D0v4BoMaYPN9C0HuyYjQlhYlp94+Xg87+IxeS7fuM+9kkHR//z4l+fxRLex
Ys2xEkm14iZ7nHj3xGCoTo7aF6Ri5FeEw549evNFSXHGoYJ1uRkIKN3Z6y9VrJVa
e7M/XK/o3Yw9XCplhSTUyHJtDWYzQSLCnNMRQV+DdU1x5KidmQOjq0tf89bw0z/1
j4y2dfnzWdzD7SkraB8X8J56/88UcXkHwaehwixzs5jHqSstkLcp321kRohQnBcC
1Cxd7pQq6beUvDtz5nr0dHH50USMsWj0fsGBlg2tvLjrJwiiCFiWX8VtHu4nWXue
btKc2rQaDYHkYleqjMg6VWrvcJzqR1VjF5eHqmEhcgAR1ggv1TIhZDZIli/KYCmI
EojApHwt4gRIp0GGZHcLAqnpUcRjYG/ZqFJPwt9a9Z4nBZWfevVoDiZ+CXFkXITI
4vQOi8UXFlH4XpaTzwfgKPawjvPNy2rj2pV6LjRa9fdjRSTngoEqxkuJnP4GrlgO
DIkul6obz79s9CFfgIoLYA59ulo5j6CbJ9KWzqyVV2zqqBLqw1ilgppmN4qDLIKp
pnBaMSVSI3sWRsL3r16ynPUBWwhxi7qutNy7RTonk1TYQEvm+vXz1xs6bQrYHKKn
oIgkRJjn9A9GrAxXvflgWn5Vl3kXHGyM/tEU3sMGmiahNBnObl3hs7k+6rrho6nV
KU2y1rNUwCC1QWk0zsLASENLuWkKXehz+yAOJ11NGBeDlUqREc/R9/KB2Qb9c1eY
4S/V1uNEaUYGEEicARSsSjAfsd2YbbMd06ZYQ4iQqcO1vQ3XBq0XDJkrQbuhK/29
7vQaQKZ7Hn0QDujbiPzhZbx2pHD7VYqk0zUkYn5Cjy4Rjar/9yr6uDaEtQPsfUc9
i4dNUWUPsmZ1KWiesBcdkLCIijtSCwueVO4HBCP8EW7TP8AAuQFi0c+0nc/P3sTK
s3PO4ZCjB33+ZdOdKUZjXfBj2F3TkkvneKi9hQH43Ek6toYPhcKrUzl0lSabSgFC
gMeWJtjSc3PyGdF43eUu9Igii90GW8AT9X6l5uB9YKPuZ0K+AaNXfYKjm79jYsfV
sKLs1naylTVQxfnOz3T7ULliz4NV43MVLpY51b9fJwcEQbRbA7cspxdJ1Yo+iHyB
KOS09Lw+1rzVVYq2PEM6fgSpztDkCujeEZudSDVgoizEuc6PmE2whb9UOKNUVqmF
u6p60xf6+gq3IvbHiwEVd8hoQQNvUDERvhanCSDVftyduFqIJkBT/g0JfN48RkN6
HtzfHM6oLcPAoTnMiiQNsK+kE7lGxv4KbB1pMTiR20vXKleBKr/u3d9ubioMuUb3
Ll1KU8wPZnIRVGU1j0MYLjGNP/aGWJ7b8eN+djJ164j/oU6Lxbuw5JZjlwbkmXx+
t7gIUp6tfOCse4y0YQxK9Tvn0MpF4h2aZIqFiQqwIt1Vf3VIWf3/JuYP1P54ET/X
jZems760jw66QXfeSaqb7QPlRmxW7LgXQ6919yXRmN1wUe1kqv4PJXF5i2nXfecw
JxqOm6XLWSLDeWK4MwBP0yvKxolnyn4hJWlwyWHm6NweQmR5LnkAfwUo/s/+5hne
22uSWDGxLNtitKX7NP3VoXJ+kBgGBKlQQQnfFIgot+gO44LT4E3LxvAO/nGoe7fY
MgxKJfsEd4/W0TOgJNKscpw3BjE3+7lnfJ2dPVSrDELJzSYcbJpjCJMLbD5pvVmG
t2s1r66ftbOBM4Wk9pz9UewBuFyoAIFTSDKqxfqZIOXj7Q7fLkDNmuyZF2jFqrr0
6SAdO+RFoEoWh5rSyC4YcBa/8X4YoK8Uh/hijA6jAztEG5ntIT4skMjAwET3AVuk
9ifF4mlK2i+hluVzigWneeppGTq4ot907VOOIrMPsN6ThuGkDA0J//eCyOMgbpvc
lr0F9+Rgh0gk8zCha8w5UgeWFE4uiiHeQ05r10mzhADoqU73k2M4JgQJIgaprfbS
YwCJqP3+We2/FFQyLM64CZB0HFKN0SHC5f6fWlUGuY4PP505xf72+D4XZLX9ct0p
r/HOzJpChqrSmEmNRMmdnvbp6qkGvy/ghxm7BIHjzjVqVYqOPqBOfPGocGfYL2oj
MkLV/QvHx4YqMQbaklL7r4/oUemKdS3UBCoRTYpZJB9d3dbEpCDSxiL/iOIpwawK
3Nu02stac7UEFCYDt95xhbv/WEXSuPCIa+ZAcPa0vPK70D9vCsb4BlMfxHJRwVz1
cR4EuMpNmw14p6s/ewnQ8nquWhTDuCp1hsGysFyIEevu/ED8f2Xb/fm/JX5zEpnn
vXgEylBNc4T/+W4hcGZ70tq0U6gTbIAx5Zrgw7dI1pShWJtXkdPexCssB23BrnMZ
L55JKmfh9CWvZEuZbDURo/8BDxMqfUBBlcVlI7NomdJWpkTOqFInve0TkqqBZgU3
8Zk2/lRFs29Z7eY7RcDRStBwgN18C2+A5bWjbIrk+3+M2xM7Fmqq0y8pw5jVCRnE
P/Iv4208rYhAWrU1MSnifjiR9Fkkj9u54xJ74yLNkygk2Wv8ORcUO6pofnBz7MQg
pT7Wg3wEa23vcydE24gGXIreRoEdANua0hj/VTwo4TxHXNXN9L9inYd45rvU3Ynz
gZLN0PJ+K+Fp/ApN5DO8Mduuk2JzgiAee7xMiZpmFMMDnN65XdS+9VpkoOP7bhSD
T21by4jo5r8tz35eiwltqDYLrytCaS1y5LmwLYj6wOebecbDmhEztq5P8N9EkTGX
Ipq0i7dUA/km16AeSY6Vss65F0zYB36g61hWjcAhmpEcL/abMeVPBJzpOgz0PiG6
siuMaaqu9yUEm5PvS/ybZLw3w+WI+6t/R6kyYDyBY13kHIYCwCUISeD+HIGvvLKJ
UZQqVW90UfyiI4TrhdtPwZXWli2pMNA3A1sYKsgtib/nqwkYkBSzx+y9v57ZFPuP
vWj8u9rsODKNsADVVNmd3JZAln5Bow6iDgfL8QcipYb/jzYbcg6kA/01HwgHUiPU
dQdQcdMzVc0tEp32pBUWRbmkVGOVlcqetJQGw52ubsMlYHwb2ju57kcjCWEdmx8V
ttN8wkd2xCjnJXs2mBs2gepkUHPFIoFIrjFT15C35EL4UNI4is2X3NTFSCedC4kD
i99MQQOxkJ9wLesOv5//DeMPjUvC5+clK5QrY0+hlvDBpkGAvK2hGhFKXyAfy08E
NE4F1aUJPcbH80zAOgHgYb7Fcrd/tnjrdSaZQ18X5s21XNLzdA+b+Y/YB+fvPKU3
1tFav4cGhKzzwa9vsrK7TN3tTOapWDPEtrzcIoAECVf+eGcDQiTGFcGaNXI3Vbts
BU6uY3OjPWlSCVhp1H22QZNiC1Ja3/w3xJ5fyXHRU4XR55KjNOhvrqcJr6dzGqMO
Xnj+M70KZLgOyAY4nAjZeLQdIjYBOCxlVQf0BLC7RTDhsJHUpprSG0sRJFXPotJ2
X4u+QaiQ6lFvODPosb7oAf19nRlo6i9NJt/lyV6TdVtmZlkz5eYH8Gw1tLAj3WcQ
17Fo8Htef93w3Zp5AjwyF9HRHszWDTlICtXCcl9gZejd2uny0TU6VefJ6/tWjEjo
AJzAnPgZR4Of5ZFDAeMqAauYexDc4l3K+4WrQrwh8o9uy0Txp+wNrbq/thiLtFcd
ypGgS7ckfAzjQpjpHZXtGzUJEG3B2OmsB6ACBeRr/yy2elmdFuauNCUH5s8YZFPt
6XVNH1Fm/+DtyDiH/Y5ByGmS3YIcjAWKLzA/wk2dWUCSz61XPISo2hJmtmxuaWsb
bMGOsNQJ/CcKRhGnuIsqnmhSLg5ePKa4ISs/Xsr4hy2wn+Lx9I8qvuSNLLWktCNU
qLF7e4j47vW2twseJ9YR+jeFsr+AXqrd4xHl7MghTVZSjYN8Cvk/9HpSrK0sr2wb
TjVOEW3rHEguArMrJmv0mE9vJjaUVW9KTkG88GQXsXlv4uAE8qXvJc9IAeF8BgPo
7xkQvn4XKldPIw+sDRUl8gks8tt0EPZ4mX8IxabRjOEFGPdJPaDOdxHyuaiBzisr
StJ+17FCaoSCm2Kyl3LmIfe67DmQgFxqCHfLtUn2S09RJJXpKvXNDGdWli1fOqjl
3HA5FGXqsdxx0ygwLEYtskUE6a8iS84HpXL9tOiIW2pwU0OLpotbfDPNHXKw4ltN
yUAolwrUXvXVah/NIfjSfdWVnZgSu+OJ7VpRrxBpJWm5+zi/kzLGkec5OMcZv7yK
hbI021yAogkiLGZdCWpKzO0Whw7oHHijFItb4LpLAMowF4sdPQKGka7U+McTNeTe
RJ9AwZyjm/ffuv2L+so2NwdBZrns6qpFdIqrvo40qu+PrbuxrRT+1qtioT786ZAV
5AFXmj6ztNqTLlypTzXlBTff02/WOs5lBYLfiSURo5l12oTn0ZCRT+K6RhTT0HtP
Ek2b08boGe9zyCWOSdQJagDZi21FKBJsHRyPldHiS65OBl+92/qn5dPVQOevtTT8
tEE/A1g7m/Tr8EOvIqOyKl8zqfMNgS3iSdGL5N4AxqtvptnJX4dDNjOx+Bfw3SDv
aAKPLi0k3IXLnaD3UXSVnorK+8XdTSg269AaWutqaultpS/8/Kgi2VEQpFf0OIYn
jWQY9cKSc/q5quSi2Be25AoP8N79z38selgOet1faWlXfN3DWHT2Vi1gLLBleMsT
ZuaN2w9rOoyQbHMLlw75jSrNe6Q5if0FXqndSo3sIpS2DDPweFQ+Mn6eNMQH9smv
DhvUTmi7grucG6LfMXQRru1KH6efsFz6W8JXYMrhBzRYyFcyvHrXvWZEJ+VYr7bq
9q4QSyqsJJlSUfA+KQGa5gZSYzxF6+VCZGyjwtIcXgtKCGgrq9y1jDJ56FYJo8dl
c4YPCrYQuFQfQxPU0hCaMY31kFEJ1nUUXnwTSt8FyR/taaBCYoskRZs9m0smMfBl
s9KXn27XOMpPHcfOQG6fo4GD8Z/WFJwp2smGZGDEMlwd5GJadkzgBptcDDT8coVw
ESG5hy0j3KfpKYg4oRx3ucN+irwJgT7R0ZeaRQjm4i0JzvJpS3DupfNYInTADvR3
DXOYEGg7+4vcNfcvzoSifGZtC4A642kw0HTLlk5NAEqyrNpx0zAe2c0M3fTLq6aG
3kPbh3PRXy5e+GFuY/apDYWIoj8sLn1YmCemmoxY6d0S2pLjZuMOKymwwAhEuLQ9
O8JIbKvuEIvFJykygfSspx/Qxb0VAkdCdwCUxfu6kZlaLoW9sCPUIRO+MWtlf5om
lhT3soLq+wBgJkUZWmrssta0KMVOcUTssDn3PmVr1JDBYk11z9S5OnYV7ReZs4Y4
jJ529kqfY0PRJqrzWvxhwayTJU8dP5ZB4aYrSch8/FeUDZ2J0LoKCSwlFY1ncIR6
wrvvK0LQKu0e7Ju84MUbF2aJ5WWM1xGuMcxMTLuMyz01p74GIliwcJALItml+5jd
Ur1IpG8Z1QJPQNsqAUqVrZFRLv4KOR62oNcfq8CaVDsM9nWQLLlBHzUXelo3jWZm
lxyj3Evs/W387X83F8ZxtlItAyaR2adp4FSvW58LlxCq/fSfSNjxjhe6lzQcjXfV
ZT0gDVj86vPnR62UQ99+XXYXd4oy+X0WBRJQln+fSPbhLGV4MspxADBxFFXStCtt
YQDpX7VlLuOPVeFlTGMt4IHMvnv8YnYfKibroOTGqr/KmtHAZ8ChJXDFCWwLLbRQ
4wqyGgWCwHX/4VVMOeLgrB4xRYSG8i58+GRgMzC67IUrnpZ2bsX3f9fsYS7XkI5G
d4rnF5LapmeXf/xLI+cR2aDHsQR+TIm8kDKAzCVgvQ/5iZ4uf7vS1strlTmpKVwN
T0OGB3KRgo9c6eiQold+FGA3EjDWIhq2VlyEcZfai6sibkxAVPK2/KCyOekg8Mof
WNt7iU4d+jJxjzbcrRQXZHNaWWghAWEqXA2aFkw4j0CfvSIVjiQCJUERmzA2Qt4X
IHrMmLHUqNo4CmSfwSQblkmGUyT1ufkx3Q3pjNMCI+YKpfqyZ9e+iCUWdf1KRGuO
lioCxDsdlI+NRltCJxK3Na8/ENJisyRzn5tRjNZGZP8X/m6oRhDcc2RaM5Ll3uU8
iEBmmJP09v4tLQTHbhwSKPT3cZJfzsvLn6K/LNv67zTpBPp3SSzoCr6DBnA6s+Bk
nhEjCpRXfuNH3Ek2oQUNXIfEmh1yptMRzEtkh26mUnoEclyagRqRWjCZBZvYoGE4
mfcVPAg/ZeCCrqSsSbJAfO2cCCbCX39y7xXYOeup1I8xPmFGA9g4ZT8xbNb7RoT1
D3Cm37frDFz2SEF/E7r1kFDugP5n5txnZE7SPS1i7emghInWf30Vh1L2UfBIx0Ri
t3ipATvFP3JkLPoj6F8evj6zu0oaIiITXRL6ci+NbvBHG8tC05k1wC1EJWzN37jJ
QNI3aF2R4FrDD8QFRg2mgteZ3uAZ8qFgWmv0+iiJDGVklGlYbA3NfIZLphAcN9c1
EQfSleSjSVm7F7RORh+jVOuembixnviQd7fwrPhs3NVeX3Fum2cjL6wTW8prQgbb
+9Ouv0zi0WBknQNwnvCrSmS7PTLuvjaYz2SOIybIh6Z6UDLULfI8WcIGqXTQRDtC
NsijA+NE6Yn32IEJOSSkvaI18PtG2V3o+ljK1H8BCvADNe5W9edxPg4Itn3XVgBT
ZdS9SY/lwUJY3/wM22//XchYPJcW7HBCOAI/JBRWkGBhvar/oEcpS/4cqdzqAX3n
Tf2TiLcAmBw45+gQohkxjB/lRLN2f8VhIcIQrTgyD0C4wpyKL9cY139koUj7HxsP
CoQ8ccn/aQ0jLc0wRn0Vor3jzR/fXl4oAvrKWm1t5iaatcgutG7vTHVJiM7LAmtI
Sfq8ZoBPnnhYXMlgUoW5LqxMXqXvbDY+r/pi9pd0o85IW8avnEw37yFkXj37f9oM
PkhI85A5oEfC6HvhQJTD0+KaTl9yIXp9qRRCMRTMNCo9n67Yj2pdB9PnnB43Gve9
KHIZTGevEFuEBwZUqm7VkNdfAyzgihVUf7vY+4YcboaHsgowO8fYEF/C7myQWhDK
PEUVhFpOKD038Iy4AHs9z1vENphjz9+6sc1Jw9oCTQMeqEQEcnYiUamQXRt6klMc
gfSlFA/3iZ95xeUubBb7R1njsSJ3Vycx0Me8tFBK+hkIazPL57+oadZiixfL6SYU
GiRd1APpp6LuhB0l32HwyjjSFhW75CbfxCkyslhurOosuCmIPLgLPeU5YlxbT9X3
egb/CShUvp9/JURw8hMmhOwHcF5l0OlAN5z2cjzfg4TCu7sTu0Olpmi0W1suTGAF
FGREcpz1hShxK4fATNJSVbTg1J7v2arIXrzziCTkIBBfXSvZr/+yT9WbzYPXUcFw
sVNDySKKha2IFM9AzD4VheMqaVv5Gukj7fugakVx2cAHE6FaeiesWte0x70amJ5Q
g7he7y3H4pRvXlupjvDMWUwu60vr/hh8WPGrOuPGDDistIdCbqT/g7c04rIY2mL/
JmYSaslKDy1VZktP3r4gZWoAtPDgyGbwshb7W0SWP6qpisPzbIUxia4/VnPbADYN
lSEEDQmz2lFiBAARBtOigHf9DxENrbbLBtV5DfRgtk3+fKFL4RfsBHlKxxT9YdYS
mLCDZQE0cYcr9UnfZkEbTrCJDMDspixhRKKMUSK3B1NRvrrSxQARDoQKFw0V1ksO
iDELw8X+u7wlJ1i1RUUeCSXK1vXqrRp38HcpsvORnULSk5GONyVL5seQIpF5cWwV
QV+WYqHWy5qknz4cS1h7BiqVK0bEAQA1v7EOWkvlV+wfEke5UdNNKaqY0OlFUHME
SNWAfGdOMRARY+1+NzMyEhBP+6ZJebcc84q2LN6pNzBvtNagZJVx4oL0jSBr0A8q
T3qtZ+qcuNj6Q7ZBLL6ffyP2HPZK6ktH6PrjzPI0kT5qhDac7N65kNDZNpAfrmtR
DYO7tIoD0PmlQrV7GX4DQIZF43PAJEA7YgUk3P/WLsvVd+mA3cDqyOtmZbctW5WZ
3fa0e8mWQdyrmywbv2pnQO9xz7H8Ug5BiWu0VuQ4sr+k0tJeOELOJjP+XOGQ5BO8
YJqDgq7g1vaStNNMa8HQEnsrBHpLTv0GYg2HJXC9qBOqMwWhJLjDvcg09jmN4Ux0
jciHk/Sj5Ov2+AJC4O5K4Vj2blEwHGkL9gB5IJheWV36VheCcmK9c2Dd0jDmmlnj
8+FJCEaf1Y7A0E3rqzAQ04qgE0oYHgK/P0csKsGID9patqT3ijhc8k5jBcN8ISZ6
HKj8N3o47+kp+GD5ApDz/aeY0LaLzFRvvvEZIGnJ1hWnyPY40qj+n+QDFI3qcevZ
PGiEgCUlMC0NGvGs+LIYxwYQjf8LlrRRRafbjV0TZDoUmZ/LBVfOa9SxMe+eVNW3
VqvsdhHSl6rRfolcQs4UrmNR3/xuPVbTbI5G9aULJhdkIRLPvffeasTTG2uI/bAP
VAVg/9Cop22v3iljZSrfeEsqdbR1h+1o8jF+X5/9JRfPZLs7ZaoJfheaknAsVMTH
7TmOkqSAe4QpBur8y8JNlVk7McZ4NBOc5PTDnNMfkaQHYgF6VweSd8er58+A2nsy
6Pleim69GK7cfPY+QHg6HXuldmQZ2oFeT/uKTscrP+DmNUAsmCJNQ+WEc3YVBRW7
5CKo5aFVswdIBrHBu5gznT2cbhHHiA618NcpE0LR74SJ+OsTWew314LnSzDm1vIj
dHnTgVk2VJ1mPLJ3eoKaQM+rSvjQtOMZx2NHf9KzU10Z/LFyrPc0bDkWxCojx8u7
`pragma protect end_protected
