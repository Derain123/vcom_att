`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="galaxsim"
`pragma protect encrypt_agent_info="https://www.x-epic.com"
`pragma protect key_keyowner="x-epic"
`pragma protect key_keyname="rsa-key1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
BKpGstnvkWMBzNzRNVzebDDwW35lIWIUdDD3svqumUKP9qow+JgWsVz0WGWk6V+g
/EO+Pkjp5Yo3D0gXGrBu8owKZ8fPz+DyrIJZ0sjSPXaRcwR9nqpOAM7xkl8VEjGh
lhY411Gopop7b2+0bYdqUi/Vb4ge3EBH91JrGR8Bx1QdlIPYe60WBq4u5pZiC3qj
gJN4eEBnD9VMHqfcra93HndqSeWI6XN2C19uaFGX6YrhNiNoDRiyF6oURagRHGNK
fDZbUxI780wW6JTtWdvxbHqBWj0AN2HXy13/DyLsfaZgB+ULiP+yxVgwx9Wn25P2
Cd0FHvVPmulXJWdS1lLLnQ==
`pragma protect key_keyowner="Xilinx"
`pragma protect key_keyname="xilinxt_2019_02"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
li8xyCEB7Y6HUpPC5LuHBhPEod9zTzKJ3OxmRgeiozlhO/HtNki+sCeABg1KsWgS
UD379P9tzIuOvZz2nVANjhA1ZzX7mo2elsj12GqSN/hV4uWyI/smjSOgGUxmz8p4
Pfa/5iMEEsYYCrJWPrpycokTl9jHapTv6zWaFkres0dJVmeF1S4Ekz1dWmxXs7zS
+KDit/FqrkeZwZhra3WKqKF1unmcYMxIAIAsptA/ndgMYKLXArIl8ANopBkI5uCl
zEOa7przGFdmhwQSGMids+r19KMtN71cyewkhhg2W+7ub//uyHZSTgUn/polwc5r
vGmnu4AyU/JCn4Hk9LGxNw==
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`pragma protect key_block
tTR9gR1J3Gl1aUIF2eKeqTwDBxKCVHfnRYoe4RTF4s9CHh9nv+7SKNp/s5Vxh/YP
KxDvtJGIPof+8VliLeaniHW50CopPNwrmOzub7C5GvTdn/DVZtUGSnlTbCxQodT9
6OXuSnDAUFYeFH0btjKMSabKvWwXiop1KXHJGqaJYGk=
`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
CLDz38PJ+UgSk58g0tqEwfOiNk0cxAOFlauOEyW0Ws8IRovm/VZlIGWAwGXscxED
SHZ1JgaFDJ7pRuyvdV4OS0bp4FgijprBH4nWSvEZI6HTRmH38nMegfyM07WWCa96
cRaIcEzDtAz3dyTQ6OSQRqRd/+5+hdG8mTvCEjTgFm1NnVxfFYiCzMY10YpgjmfH
Srz6F56IgtRZIEgoCo9AbVgygOf61UHlbNkgVVBeE51xHvKBzT2pFNnB1jAma+H2
XUWj4E1NXdWka0MODlGe3nFDnATvD5dRMt4YpOK7cvCa6EFf/smUDFOT0aWoh3W9
zF8Fs+3QGgt1M1OGAaBpcQ==
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP15_1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
udGgvJ/+dN+UZwlPo7PwzvHeF7ke7rBAk2ziRqTUMKcR7RDwTjxqQREZ0MuW2Xut
AsGz/icp6081F/CGHLgtoJsRx8TYJzSx5RinfU4XbxhC7B8dYqvwxHdeyqOXCmDV
8uvtDfLoKa1UH5sDnvfsPjR19rVzG+ZnLtvg52W1ZWRCMUmngZZ1i0BMXEitk9YT
tXE7/8swmcPWLguI5Uv8yvW/8N+P8iVtF46BCQPjSvR7IqxIo1wfmgtoLWJG4bsb
x7gSTlapdKyCKpPwuWMImgA7InlSuQBOYiQFknucmP/wJWIPG7+jE4p5/tycwfRR
FvXKa7WbJ1vKaKizovZk+Q==

`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 960)
`pragma protect data_block
4xncqfC6E7Gz0wIcw1cOexCM/CCVP3VfpP1GQSC49MN2BFNlvNIftekEm2DU6979
90D2MiXV5jRILZGddtJfrOWEV9J1ucvVZb6Zz9uVs0TTiG1zF183o4i3wRz4bB4J
UmX+CgnT4Gi67AGcWgULrFULwDXo2n8x53hOpNM1eY8ylkryIrjvErwx4DigfJPh
gepL881aCJ3tx9zB47wPOA6PSojV+7M/p/eZtHjbHcmzZSjvzjv3DmUp1dLVhyHy
WrlYaYPTnn53H26uveVr9qQAHspmCheyNWCn6oadTIBhVzQtXSterrX++T0WzuYZ
D5qChW2Li+MWY1O80peTDpguh+LeSaytpN6qzBNo+6/HW/q8EWkk81ArQyJXw+9x
6X9GoijXhWn5Oh7I/bnPuHHA3L/PMQOVhoQrorsgnUYESSE9IPLvGw+eM183W8Uj
RtLMXKh5qABJmCsbXcfm/4s0SwviQsUAPDgVXNJrgQ01nsqbFSSnRm7INmS3aUh6
t4tA2IcoFeP14Pk5YoXagVxGffEyABDf7d2U770mGjGAJcU7ULkDZqPQw9kkk7Ih
g0mPTU2dGm/+9jqJ3Ed/p2iQDnzmoka8GcD2a1USVIyy7/YDKDuGzGIc4m1tgp1l
TLggIUh9WGtNC7uuJuLEP9/A2jrLpkcDCM37mOaSUz6aOOfeQ+QJFp3LXc/L+s+q
/h61SklPFclc1+fZCc+wJfXJ0zddO01s0+hVAA9Hk+2Q37gCjxh0ZGT1RP/+bmc2
2lJORbr7NSABqAjYHQv6lsdDSGyGikj4kvF6bTfEz2JNCxJIn6/R9wIjGCYr7iUh
1l7EAsUHyxFr9dfubKiXD8545zrc8cBCSQrM2IMk7HyNvp+N8TugLkvsbt/FA5pX
zuZSUyBoYR7CZPcGpvtu4EcSq5wnMEU6I2q6QSLpK4kEMon5ZQGt7IkJTeF/5Fc8
XjI0Rxe7rCtkdzdBUdFlCgXL5h/7WUw2ZsH3ANNn8STiiZv4fa/GSAU0DY7DE1YW
P1XNfaVMQudvbqzLHIcu2Gv2pnQ6TGa9v49knmIlVPWbuVEJNjSF0Mz9wTLeOLJp
FqGqj/8EdRzj4MohT8nPvPOVCCqvFkkSOtZ7xqlaw0tFK1HL3GP+T4Zh8+dM03p3
ZPPRi0qHm6bqh6EtsY9v/d3WGY/xSSQm4SLC0xN5+6mQ3nm7piYcFtO4q0Pb1u0R
YUnTyhNohf12A7Q9RXS2jJ4GrM81eZ4OypA8t9KrYl36i9l2wj32jMNhYc5cTPdr
`pragma protect end_protected
