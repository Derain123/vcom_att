`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="galaxsim"
`pragma protect encrypt_agent_info="https://www.x-epic.com"
`pragma protect key_keyowner="x-epic"
`pragma protect key_keyname="rsa-key1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
dYDzj9yiyAWCOQXoP9INljESxoo2Ch9LBytPTRoEGB6wCTU4hiJH25Q4USEyTxoc
j9ZPmmh4v0Jl3U2sECMp2yg3Ti/ea6klhgwww4Q3KKs0r7qocel9QBJPibgm/sHD
r954yDXL3LC5Sw5nac0zsWXbgKVbcM81KKHL4ON7gQoXzSRAyfuQc9FQ/tmNSLbH
M/xT/Q5cVHCU846apsFh9LGp3vQ38JZSaM2WY7XphrlliOGJfwLDdoqTS9qLLURK
iLXucQafrTt4cGUBTr7nycYigSw7ZdqHZLP6KJWNVdmxh7+INGLQ9RZzRbfj9PGx
Fh6wmMrT0c9pk7VYNwM59w==
`pragma protect key_keyowner="Xilinx"
`pragma protect key_keyname="xilinxt_2019_02"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
HbOOLBldwRBXS4hWGRYatZqFar4b9dg69gFwTGiQkDPryJZOyGO5swZJcZqIK5QP
4EIDWYMf2Q7e6VsjWlK2YksZ5ba1kT38XN54z3CRAuLZHJls8WvR/EsvgSt4Jx5Q
tKiNJ9celRGoLu9qsJAcwTcpTqOCtRbRv3Aa4NUFI/uqGBw2u7rrLF99F9iI9dJI
mQHug+0dMRvd+dqCCefAQh8O8L8UIEFMmumApiBdix8Z5LxuZEBzyN1B50m40Q0K
qpLz+G2bLGvYGhq719GqNWTMr67qC0yw8HfYPKAJNL4gCtB96Em3L2x7oemrZgw7
MhBZaFI/Zki6qH3UL0iPCQ==
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`pragma protect key_block
XLd8v0TYHKBkaIyJHT2yww0SUcTJNKjcy+F0eySNLvhNXyTNxlr5/MwiF/cF8t2M
4y2ubOhyJdFEWNg2KFsIQWJgNrUGJXIbeklNPpiKARtnCdoIG99RCXuNKchH5xHY
VR9RFf6XD8BDiUz8RJMTtHI1RK+GtCb6AvFEI2VnS4U=
`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
DcQ5VGUkSRy3mfmE4lZ9+ldYnHZ9F5nVpJ2Iu9hhNla4kT5XSyocs6DtbF4pJTa5
aBP9JE9k9s2pXsBI89r6vZJux0GlhxJPD/PEMst2difciVYezqoOLRlTFQEp08j5
09A5urLw4CWRz1OjyiKwgpLpmKgPcgItSu5ALbm9WMP8ky54YIEe7u44ydfbRR8Q
2mQoxzbGnbu0YggkpKIfZrCkWB0zKxsgIwkIJ/hNxCrjNshm0yGHM1JEi2XQyz94
3Hv79crBxhT8aBhM1KgRIfscD6YhMRN/0m69AKoiwHzcEoZ+Ltgxsrc3mYKbqm7Y
JDYReguS8138JKAPl5imlg==
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP15_1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
taZ3O0Xc2U2esNHPRJHyz3wAGN2JoW8pcbxj6Qe2Py9JwQWkiWAUBTLxYxs0geLS
7XYlqTm387GXrxvEWxHjv9TdIg7fUzT9A95le0wNlmqjnEG9zvIDQN34xvdmiD6S
qlCZ2Lsdbcz+aJAMz20RXbGAGSEoQZYgqlbIIRFieYu9LnpTr7zdn1MycxUhiCS0
to0XeW6yuPW/nXGteQLAUWdRrhLbjS374q6bduQ5MiRzejsJmTqxVwym/Nkkn06B
Wb/p8HB8V2Sgy/OM3Qc8nA40rlf8wOKb8QYeOH+W4lCA/urz2ZeJN8wHRyyYka8b
CxlOluoaKSZ6a/jwwSaLcA==

`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 1984)
`pragma protect data_block
26+iQIh3XdpeUo7R7Ctk2kRYAsSMWJ02VFy4szQllObkNXR5JTUk5yTijmKg4URC
crcAMV2T6b/wQhKV0Vj7zE4PovT8RWDRtLPXT6iZHa+aA4fIDwFFRJMgDHqZgwIh
YEG+sO7TFWvLU9/TMIMl8hpYDEWUlI428mqSezLVSt3WCxIekZ8ec7R51hGkibmz
Igfx97R2MuJtV6DtlxUtYmgv+QIdEWt6U1NbJF9ikvI6KAI2ypnCfKXiDf00tUIU
kKwQAHvPhTVXlo9nwP2wF6dgZfYpcEopcSrATjDA+REL90SYZSmYXl9I9crSbOzw
ghic+3hf89OghyoXwIxXcirjmvz0nSS0z2qhzmBffd/VdfNq2CcHKvYQ8R/1MUdN
vEoE0E5Y1rjdsgasV2h1s638sKGUptLaQmX6LEwo4KPbvfU1h/1g6mV68a3WDt1w
uAA7iEgmbyJwdL5ZFFTongkqhN//LZW5fYMBLrkB6XbJ/bnV4pX3Qpu6eSQn3oR6
ilrA7BtASEwFJGWNlPYarGhWLWgszDaaMFAFa6sewTSi4n0UhzxR+vlPXMuaFVrd
bEj/zpkkI6dk1id3zTg/1QJWOAZZzBZSry3Z4V7zL9zS+0AM4Og10ZOez6k7EVCF
Tz9zjMftDFqb3HwHa2OSWT8z233r8OsHUeXr/waC7cxMLcZeUKmeSBWpalUrtI/a
CPj99/P1Y2EOlgpj9/AUtzStv5yFQ0loWCDumhhwKSyfa7HVhiRkp/M8EIJOiZFx
WrC4cEs99naS3KNCLe8ydkaQGGVAKhubls2ajdnduEFpQZmb597iEOxE+Rzc530Z
dg6gS9i+pex+vgeO8zUA00eT6Fb8BYkXjmTdp9FfXGwUYie02edW3Fvr8D+s6j7A
HBR2Hf7AYNJvbFqEfAct+O/wQj2k0sc4LgVzo53Q1JEkKmYiNP1p59rM557yU3Pl
CW86BXdXR3MTEI1eNG3EAGo6CPpx0ITN39GEHsIgSrZaKfSsu2SP9foTc+kP/xrg
pqYdEYxCBSsutS1F7Ni8U5VMWWn5dF7G0D0DuPelx+fOx3//yOo4Hm5ZTdWLt4Is
8eBwwMp50taDIELGgKk0m22aWuXSV3Wqc2LL+Ji3hnyv/WV/9xtm8TdQ80Sww9ua
1hCaNNuGV/wawCrZAZa/u2UvkUAe/z6CwgeQ4PbgWVL34IP4A4xtPzQy5JZo69ym
dlxsZg5gWKuoipXgTALTPE7P/tLuqwqry4kMuh2wtXsOqJ2NxHfX9L+ThJmdunyG
3VlkFYOnqJGCeFu1x9ocyF7Ym/BWvGpMAHv8wXo23AakbyKJ6RYmEFiqTweGN66o
r+BP+lZECY7LG/XwiSMkQy5CfmsMOlmK6aGsYqa6GJPRyA9ni46WcBQUMfyuhnbo
6l6eRC+MrHZzVm29kev1nALNvCTBsyjGEyEn/Yzg369tVAeXzgMPPy7q7wK7kHBJ
/WyiUW88PcvrxO5WKw/lLPV1rBy2eM1b0fYkMpH/Mbg+q1OTe+I+SavQ6XPeEABk
NKBVx30Dh92HI/7EAJ8fJ/lwjN5C4tQejpu45teqGzrvWG06wl1GykqR6PrGWgwv
2ZWS0dZ2aZZxGC07n46xtN2mW3e85Q9uLudKkBF/9w0VJVceeqGXYLP7AOZyVo41
EKH5pT5Mtb7sv7ZRMPwXbcCET3US9sqM0PZ+8PXyn/+zHksozLre7V7wEWqZy99l
PJoXhrkvaMcCGYxlA54nfNY21imvPa2kdiGq6BdyEK/X21WCLeV8LNBPjHs7gnTb
mMaIRMgVJks+zA8rEjeB7ExGKUJ9KrEC1ssjdga/9t6yB7dOJZLWNkDhRBE99qHS
3+711B+B5kTXe04sI+va47gndyAaOnWAigeqtvMa0juwxTvdy1cdXNB+Q441iBOO
FnHSvCOQsxZrSqjgUAwW6Ds9cHmN1nocH/7pMrdnKv2n6wMColyJjWYVF+iJeowq
pdW1pQhAQkSU393yCrdsGs1VRwbjqpdXbyXaAwvNAa0mBDOWYueFWZYzF9dsfV46
IsGEBk4dBjNrk1rikFoLsTkbaQ2rHATjFSK0ceIdDqyCthcerymp22etfXZJcARU
ik5jHONr/oDJJ5wQKoirzmu0sgJ07nAUIrV2eQJWxYmYinSyXvcSZa//GPIeb1VY
StC9N1JBWm723b7c1EQzPDj9j+Y+TYIIboBHo2mhk5hKfs3MSesp0V23+nLGJLNB
WBOprHjb/AW3FGRdW8brPa2UCcsfNfmcSzaQFx3g4SJxhvcv703i41lxoe5pwnPV
lJxOPejNcrbspwS6IkSr1jghTVvadirEnAXgizRjh6ugGT7/0pEsmXZ03/NQti7N
skqyd5P2a0pITbnu9e60cMKPFcu/ARHAV/qT5J+hkb1YtpRAVwWVSbPsYZtliDlu
0+GZ3fk5SNRdp5HZK7iNn4doSfs2dl8yd8r/fsevNdsoJyg7BxXapI0SIpf8pskw
YcAbmNqlUYMZjmCOtIagI6GZXvbagK8IzjNns+ilflloGgqF0YOElz+L/19H4UZw
aO9NEdfXpsfEeKPNBOin201eLaeTDgLFH+Pw7eL8c7CtKeQvaka3nIyGbF1Tv2Sg
ZsFZMmxewcoPagtDSa7GyA==
`pragma protect end_protected
