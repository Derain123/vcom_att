`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="galaxsim"
`pragma protect encrypt_agent_info="https://www.x-epic.com"
`pragma protect key_keyowner="x-epic"
`pragma protect key_keyname="rsa-key1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
ayrcL9r4O/THx6JPP0dgz8L7PylfdK5wdrxfoPXFC3ByY/Okr4V8/6IlU5+DPYY8
iLf7qofEV9GwRGA4EYPzeQAD+NUkZKfwWGt2W3MdZQWLNamaMfSH6fUMXedewOWf
PhM/qaG+lHO0LSOCtEe1mdRoFrvET7QeVARgn9+oArJSu99SG8J2zOH1C6KYKD3Z
BmE67f9tff/XxD2Dv60MIueh0nUdAUiOarCmg8lLRY9X72rHNrJYX+tSOVtFJlev
dLt8pHIenAbH5PjHlKBagz0lOLwcUXmstzMeQVoRp/707aY1DXi+9xQvqcP+D07e
OlGkITHSP7ZGwL3ModQoSw==
`pragma protect key_keyowner="Xilinx"
`pragma protect key_keyname="xilinxt_2019_02"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
QF2J//1k6j9WUGplhLI8SwYA/+b6RC/WVCCU8QKcKuyB3f+n+zjRsw+KLXa6gQfW
gYiNKXdOvKYUwqx2tH7fR72vSeG10YQBh0x9Zd3NtJ7GQIBcJmCLLTErVfo7uYs+
asSgajLG9zhETplHR/I3RugOkVlPuUPLGrBSrfDmfodYFaoAu9iA4TXRBYlWSGOg
9aKds9BSL314d8hQrFcw67UnJWP5xOIlFcrwb99Gr4ACAAeORcQC526SPvz4C5Sg
vN2UQtJm2r2q6L6ZyVbEykbxiZ2HUEAMpcLcmhCgJ8JvyRcZ5pENgEi6N9LBiMqw
kJQNuQCDrCM0pF9AxJ7kqA==
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`pragma protect key_block
pNCzGHi03cWreeq1MvE5o+YFQ2L8kb2R3ju5cJbotDuEasDbsfAPe7Y3nvzmlYdQ
eawbn5i8JbQH03vbHTCUV0W+SO53Nk2xBQLh1kwwG6JQvPZqogljJGY6/SDh8Glb
nm+tPi7l+xZnj3PQgzdH9EPVhdcmgCYKLldqGk3ZDtY=
`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
RffjjWnsljtfvX6LCVsh69V7tCUXpFsUpo1q17u9YIHyMRy/WOHqFCUc1MmWEwaW
Mc8QmCVLDnVwRTFJ7+QTSCeFfkKXxR+X1uImztIUcgOEWj2+jJzhdRqeKzaUOLFQ
kqolM1fJzF85JhZa+ufLo9mSZ2vcqKaQ/eDX5aiiIvb9KKiXDYit+c/JxoXUkCvY
iNo51eytjAl7roNqadhj+BpbQgVKQkVd1SxiYHkeAI949b4y60PLZXHt5IVVPDEb
8TjBTaHbg60Md+qcYJZvocoRtfxMyiUfgooQPhwB8gYbb81XNevJra1nJ3cfjdrp
Sq8EU4DmvuZM9a4LQrhkxA==
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP15_1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
K3mmzSrhVpkh5zhbiUaJN4HKaib2HWThmo39TsmofOHiqf62V+QLZjoJQrWexCVK
SUBmfdZyvZskb/q7d8iRv3R10deZoxx+ZowRfsu0Yezj68lrNNIJ5X3jPfL/TTsm
0EzsH/9LQtmGS0Rgn1nyZ/9C6XzGGPoUstKvfpY2sTWOJc3B3XJeRX8XkZoiNK0m
hXb2glhZp8tCNMmrrPegLGKkRpqdz6Ln4kSRHdhtPHJHOD9swD2LC0eNsTRoqxoz
jgn+p0FM96sofeTUM7AzE+Qw1+sniAH/78znwILR2aqvxKJonZKVz3MrAjXQ6084
MLrjQ53xwUFibiVOO9FYnw==

`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 17456)
`pragma protect data_block
HFIkxJCrRaVY23s/kK3fEvrU8W2ZRiZBgayQQhdFJ5/hPQz4y091tw8aAZRfMjtN
Ed0Lwytpow85Hlf+W1SGTMlN/rEsBbGHz3zd3pHxvsI6VX3HPZzlZPfpWck/Ah95
DsQipw8Nh2Q2NsjlFcg7amS6shfcb0baSb5NjQ9fdcSMGGyUUhaPRLZqDMmcBMxz
UT0wIujnwOzBwqoxw/ZIsYh+HqVVLvxN1a9Mlmd6Im7KV0CJL6loniIVsVNyQBdw
XyqcNtA4IqIT7dxxR8fhZA+Ca2Qkef/Uh3qdQVt+DvuB9a51aDOxHbNxZpYE88oD
/pvLH6JbSWbDaTO5hrJCzsjlEtKe9sNZrMwQxqNJj8OrJa1fYfDGScRCKx2FBLts
DBo94j0Bo5WxKmn5t+Jluuc954cyhujsE/NsH7aSY0+HhPNCv15Mw0AW9TXZsHY1
GLrtBPUV2Mb0gZm+PcOzpI7p3R8v91wD88tEuOlFlbyE2wyorKQBy8RWZPgUa73v
nVbKNzcs+A/+dhdgBnD4rLnfviYQO5r/6AnN8LaR8sjofjpwKaM7dsnsLQGkzA6b
oqMsnsDBGc7Wncw3RJsSRkQqiNfagujwyazG4KqdcYfblZYt+Jiat7dFYTVJEPGm
RGOO1Y/tHUUE1HdNhCE3mW7PMhzt79Yv+Bkl/JNcalOM1yUESE5KbUavlXS26iLV
74a4vEqK5fSRE6TPy6MMcOuteHUu1PVGDzIZIR5DK22ZD2oO6gdwq3RmGY3mgSta
UpLbUJb6Wg2HL77K1SjDqCCpT0Afmshn/V8dkbA/5Q8saF4adaqt9U5Rkc11783o
w/bm/OMzabcWkjJAutwZQxhIHIdjt56C0DXeSOlrO6InHzJ0HiSUC4s3AKlOXhVL
P3eVEZRU+INKDKM2Fb+OfKmjtVnZnzqz0UOFR6FRwYhXmqltvYOHsOyE91CJus4d
FneyxqtxeWhjfo4EyNaO0RTWfNOu3WzY8MT/i3NPtwj9SICSWK3KdV/wtipTEfD5
7ApxeI2Q6SoBFaTZbQJ+Ql9sDNQMFZDHqxeJHY3otpj7QtbPwxDoqSZm4L4BYRjE
Aoeafkcev8ind//KJQejZMV/u/fhtdchCWPGGWigKq2WV2aWzYrEp35wmKjF8Qaa
NyWoFFexq5eVd2Y5gdLxzwJ3WONeTB6wn7GiMMQWHGAEVKWtZoCylUL2fFVoIPZU
2IWUaCoxiZKB+NRQoy7xszBgCnFvUjvoMF6AodKACB1O5ceKFtSqFXFZw9Zir9y0
PYZx75mImoV0wKOhnb6eXNbrHoE/YrpUIsySzZjsL61uneXdTrhF+48SfQPMS6l7
n+aOEVGHQhVz80mcxcOelBrNMGf4Tjnws02A8C4yWETVhss6jNbTOQuwUq4zYDEM
NqJqyvSQEwF4hVfIKepMNQDinoDm/K3KBxlXCntMMP/HDQYJsjEAZRwiI4w6Z1g0
vibfiEhWiIyJIseQWJbxBxPEj0UIHd10JVFr81UTBr8CpxNBwutlul3k00RupJv7
rJw0HqxMjk6kiNbAwyoziQQr/yq7YeP2oeoc4W3m7ZQS6Lnc9R80sMkSVZbGrT1z
E+/hk6WD/O2tgmEyDPcAWXbfWjow/oyX3uY2BDq+ain+W33/r8SWD25FH0/y0fIg
aaMxFmJgB9c7p3wTNKMJjqlrq+f1HVPcZXgxqX/oz8QX5f66PbWHpTjTa8CGZYml
Mhmzf34EEeLtWZQ1rjjAB8bRZWZuAMECGXk/piXeSS3cXh2+L0qU7uMO4fGPdmai
xzUVjaFaBa0BPMxDX8uh9/SDA8kwRASfJNEROkXk9E6VKE/IQR/ZHdJP4Ub02hYj
weE8YrLsvYxKBEOY5hRLHn6LrQtPsnVsF5PvPBUrpRVubPkxHUhvSgNa45DnTwXF
Ns2fhGCXfEslsnigfHZ9efUk0/H/OVmQXt/z66M20t+3Iy+giWTIB1FYbAJpHT44
rHPKidqGer9L6TWYe13iaRzJmIx9vzogs/cqzFfMG6z/8fz1TmQlybCKkkl6Lg2q
BEF54h1uw5VYgSDhA0mEMNBUBPxurt9JVte9IbOt6h5Q42x7D8wLQ+/rFOOCuoQ2
0Z6w8cc4cSJOYgerJCV18L+HuIn2rXhWdb0mQXBn6Fy/z8i1HxyInbZ9rLYsHGfy
M8Y224vQxcpMvaPkuE5kx8bJxadEJewzwK3/qtJZf4xh4I+SLPRNc7lyngOtv0qB
BYo3aqBrpyYU/dNdTib6prbZ3BxSvz1oikpnI7RjKU5lrFI3r+UES11ko7P5oC2H
69bBSlbS6lK+11pO4bsvHnIFDGwUh9gpBsWQT9fyd8/L9KTMbWVMPXUN4I9btp3t
4xhRaJu4gZzlspm3YNtrNQNzV6v0FDae8Y9YD3dDJaye6pff1RtunZPvpuZmsj03
hFiA4qwwRu0Q5vhfhv8v0R/XmQm8gJ14tA9RqVlhyMThmoisdMTYS0BFNBnYTzT/
LVkPaQKXZlQcFfygexxHI4WtiS+EeQtjtRvH8U56R+2O1/1d1XtGeqWNujcdbryQ
st5u6jTZ5oo3/oozmQuFVAO3EFEuEUIkcgvestNrlSug2FY9FzSIlBVt/LtvWkxv
knFFyjwuatfQoZJUz1ipXTeIPt351vW8O0m2ODUnEbWz2HjOuZc8a96SGlVzQ19E
liPXW+OitCl/JQlUZZuWBx/xOONvvMys1AfqjOLzh6RO2/MiM+o8qUaVkxf2b2/t
+WeyxemqCkueLy4Ew2GB85GjYW+I2MjOmh+TqL7dYjpwANuA9i5h47ZalPAc7oMD
Qg5Egiz6wbD4nyMxh/sEJY5WZzokbqt5t4EqGtbU1MatLwWhUgtEWyiOf0e7Mng5
E0jaAT32EHwWl6CzJCTZL0+JOLH5Zlzl9yPiwUN2nseDJTVhmhza6Z7aRi1SNXQN
eMhW1RXtGp8LLT4g/uyDxsSNASvXWW4M5IbZaWQjpNJCXlZHx+YPP6lD409esVL4
ZTqP0t02ygLaKgasRgav6SyIAYACfP3waeoU3Zp7adpJEllrnLwUnC0MhCwpnpsc
+NhXeIVjxO2drYA4r9fB1c7qkU/JCdO6XU5jLz05qQdJnnOMHWjpdputmdFageBK
z4u0ieGj6kAT0ip6MGbzSTTXDVkqpEFAb7XBSisRaTHoFm7yXf3T29W9D5WJoYZ9
PDrPQGwh/v0oeQmKYFfGlO8U1/thM51ufazWysMYeQYjEuVsTczJNrhi+Uh8GHdv
1MQnBpRubGTeQwsp8vjEU9Opqxd0Sma8P0mNR7GAOAzp1KJrzO2TsmJpv6zJ1xmk
gnTCnFGe48v8qWhvibyfeSZyuSIUaIm1PxtQx0bczfM3gAPW1fef5zVctgWEXwbo
2WLMblO4cXOo7YloklmgQs1tdpXOAiwXhjm8OR81/BwNLokHcHoUjzeqP2IcGrwx
LRD+XvoPwbcUaZOrIdGGWutukfyiQbI3gDVwpgQ0KJtztAVXD7PNPNsVzY0zoRyA
YYqzEWOBM3bcuQAi2TW0C9/ugwXk1rZbo4Qq2VttAqxv36psWt4E339PAGhs0V2j
h/Y/h1lvEr8qAoRhlEZ5cJ8Mf8Q9DxiJvb1QuWzi7H2zAXByPgflCDNT2D3TY651
mr5LBJU9drvVHNS6qQ12TDNNYmMntV+ARfhxLyhmxL9QQkSnZkXA8GV7fGjC4P/f
NW13aUli+dSIj6JOFgG/+Fw3cg6+9cWDkPsIxGOgG15XiZnnlPSGhS0RieG+jARK
+dBd+Ii8ivZ0wI2Q8LfY/sQ9L+SzgFUXtfN0UdNNU7T9oBvdpvIbSEUc4TcwZ8Rd
T5mkZJnIM4XAmnrcae5Lz2lHlrmVbs33HS1ZX5dGLMFhktv2fkE6KKMF+ENcHa7y
nvXi+Re79NirYu57Q0wLKHvpmr9pkia862zCttQVvZMBZvvLHeXE+0HgTmqsIg6v
jCb/T6iq8zuyCNbCOzqiI5ffcvjHkRQ4WlHBh4oy611P7xLgifzDgIpDAUNatSJC
i8vFzu82SMbJm8frLL3uP74A52qzTHaLT/0/jhYzqQ2uOTaFFRbL9GURQ+FpMPen
G+VpTdXO3vh+qKZ77FJWHhRpnGBzQtbOjdO+TvK+WWkgHxGD255FqM5f/tK9DMnt
UF7p+An9RVAX0d4mszsrPTF/cppDG3Ciw0Gsa27KB4QlN2EPzYWAaVTB1zazUXAp
Sv8/0dwid5LSo7d8JIMlMnzCfXNhuS5NmjJQSOWdMzX/zE/JRmyPkIgyBH0M8Fox
pDkauWhneRXtbgtGFOoOYiXUJy8IoiIB7o/Es3+DO+NslRfeSRfLzQTWG35r3VA/
bAyHrfrabVdvxrbcviSTi2+Y89XFFBLbTuKF3I70WwuEt23MAFUZjGQ3PciV17nw
cgcH2FSZS+4eJDxM4L7ptEgct2GpJM5wIFGzwAKqUNroodLlV20i9xTkCaanpiZV
u0Vxlrh5FOl7bPTUPXIwM5Fy8oSWmxMtnuQy4k9WiCQocBLqMdVpA1j/g+vpWzeS
EQhV+7NL45d7oEo9rIDiDeRvk0ORcbw/L8kPK/gljITJw9Y4aSQqBLvIgBysiwxB
tx2C6nBWPNVUrGFqXwZWwnlI6t7/a4xgTKOhEM2v6vMABp9JG6Jccc68KGillqap
xIIox+e7Daw7QRYsd6knbTq8Q5YjtOJ99trC4ZJSn68b8yBFOp9J0szWuNdv6/LD
L4aWqf5ZLBQ6mc1qOfcmH93HXTPzVJ0e6V/5/slyZgi12a8BhuCEQI24kg+XDWuB
boOdoY9Mg87lC8a3oOgKeBd5NfMJUd7dijKCDT9kJ+s/Bd91s8F2KM2XXsj+5wxR
IO242f8NgsXBQBDgYR9gGtm7ChlGq9qw93i4/m/L9m00zas69TgY5jlOrkINuPk9
6UNW/a8RF+CksJsQJMy4810/MzDpb4demh8P7QqqsxwwprNZerRy6Fk/p1UzQ9Xh
4dMTVC0126EsirZ2H8XV8DwAnskkO0n2AQfC6nz/KT3cAvh/h4pfaAUath/mq9MF
rkmaWDrfoaKO7k+GWaoBCecbxoeKGXm3UE4htlR4m0mBhrImbZUTHwBpog63KaBo
rZOatrr54QOJMpdA2E4o0cQTCKDGi3fUHx+aJxAg95UM4fIK1YVDPz2NY8q2qUX2
cEPdkcarwOiJsrG6RPehqhl9K/0qdQCSiV8vWhBIvYvMSNvt+GLY0nT1Rm2sSccl
htF/YC7AG6CTgBU0/awsKkPa8JL/O0S0A89uRLDT/+4UJDDHzXh96euBEHgytJ6m
OPwG1yZoe3l7m4ov1CEOoRy2y9zGeoOAHKTCukeVCPflJ1HbN22HB5Nurdl7dYQB
HpYLI606xANpZqPyC+q4wSYfVeLzMflHtgFO0+Efw8/DdMnyX5F0TyCFvx/LF+ct
gRaUwbd2DaRX9c667wV2HET2/nZZYZk+MrvD8SicV/uw34nR/zNhsAcNo7969qqY
/7ATetVj9jycHbhdZTsoTDmimFTTtsHB2WzyWNY75uQzSAZb2jspuDjJON8Dcjnp
1ME1WlSD3NhmXBM1570mx6UuSc/cx/d/600ZHrYQB2C/2x8eNSnLAi4AAygfvOCl
1xydws0077+GncJZJWvuXSkTD1p2XjI+aw8DjFVG+BS/pBkewdyHk9EcdzHMVp2U
/Le78/tRtI3dnrxiUvxDtG4VSO6zFALUIbMmXeJuszyijHcIbu2CQlQBQmCbKh1n
iYrDfGnhJ2xmO0FsTZwKmJWdPr4Mr5rJR9cp9AtM+i1lKRyjox8YNfkXaq3B9lc1
OoqYtPsdgJqiUXoK/7LMoNxCbtmkjPQ/ur5IH25ET+tE0yIc8Zm34MQymofG7rkG
8egqJBe0t9DyepJogDNxVBTIepHb6O51+rosfplzr8lrXK2Wr00UKV34xM6L57BK
vNARaNpint4QBQzy8/JnYU8C8yMiUlHB0+nW2c78NaL89ebygBypP5UpyDkEdJEm
+zs0ehwK+FEcLCJtHvdVtpFbPJ7W1voKUTX00gACiHRmqunGF//pRlkNz0Y0PsmB
UhztwWnSEwmzkpZoHRfMzOds29CE5ILrKK/2CzGKdFyYYEN5LydPygd87DMgNxy8
wK0xzYChM9YapMONP3PEVathLLVd0Y4Yh6uKU8qe7KZx8PYQmEXiXnqDhXYmcIC+
1nftkVUzLC2U0Ym3fGHq7zZinB5GGJIsWDdRpFoFQHY9yNSu3THOdm57eQIaJ12d
iuaXBMQBxW1d/OQ7GMbxerAS8a+1mse5JM/Mz52wtdB6nRPK1ZmPlK7KWX5wbvDE
xVrcX3D/yk9dzIr85xGIf7GXmjHJrTguQDjNzG2kUdkk3oDqUtPExr5fd7H819xU
D9MZFZjAYk++81TrDbDR66QSIzlzs9tjOHN7C/WU3KHnYUnPVjcDHCz7rddjTP7i
G/S32Zse2VnYvPxtDJtUS+ZUFeff5POngJ44vi5/jv5/UMIQ2SqfgCA1PPtvvZ28
AKsf1ke+xNG8XZuS7wpZp4ueUuZAZV3UmfKjhbuvgrZm2zPUckRKRPC332czGAzI
b6qvATfclEVCOFz8zcIoi5j2AMJSpdMLA+vGwCYILrF7xOSdHEngGhUqBezbQXuR
lyGjs9MR8uXH6fdg1YTS9VlxPXZg7/ErMXSVJrV8Fj6IvSqHQdAXsR3oSIw7vmO6
xdXiuKT/WM6LFBjq++dx3497StVeiDJ9Ba52IYppTsNXzdZYoTU+WD9wd1sG4K0B
emPq8RaM5tCrbA8a3mztqW15g2M6YVvdskq/2HoNSav45Q/yRHC6t4+O/68xK+nj
E3hWNYTDGooJPyrufgygqjzOSQJyUDV6IGOoHrptBRV99qEUkyTDdaVZe9T7VI5q
LgQHz3Z77Kn7pv0A3+PUqbyWMlSgqMRfKWn/VcNFwl9gZUFxABSS2xhN2sMdThuO
0jFg3z00Z5LkvexYCmdb43cBBa83jvHc9zRCfM36+DjRnRVgPlAjnMnqkJKJYNwz
cb1y/XZ79qpG1cNUgrTW5UFydGO35ijB+hFGZGYqNNtcMBP1N4Rnrx7tpNpzwK4M
CzqNGBC2+dyKkiD68orQ+ty48UIyDDlD2Qk9DYyY19CsvJNfzgtg+pYgnzHbRBiw
zVKly0L/CDOI4pyZ9yjg78YNfsPvv3an7rxhsEzX/hYVaUgYT7W/7MrBqc2TijQQ
sq+BRO2hwKNFRrQq5ZIpD+aPcKXRbIRiLpJsJM/gyPrlyONZuemWKDekzj51WMDZ
WcC2wtcP/BSctUfECos4EusrJ27BQSxEu1mEqgxSsn6Xj0TFEGn7kv7APywbC4G8
PntulsZZyx8FGVM99JCFEBjVUS6ZJyRYIaaA6EA8BKLxjWRB4hJhbV0bRg2d6OI7
LR2YAxcKDiWKY+R9T0VU7/lKkSd6LklOCqay99TnqkTqLTdnMQvymK1F9VgPyArj
TqNwABPyzZ45VyDjYzqQvkOwZ12qQENGzNwitM5Kfg3q0slLnVsIXvbtX1BxXm68
NFjrEPIpndyWN45NAVUHmod/FNvD18/lXrGbMoftg+IrVbQ+NbkoHZl76HkXtK71
CAnoILyDOu9JwbIOFL2uO6wBTkcnMZ82VIIIXuLXUzKyPjTRZWBLpWsAy+M4bU9x
M7M4VUuntrK0/L7249WmEBEQ7vtt25dG0FOtZLSSZvqsy71VWLIm4O54oFJ7XQLU
MqfCUBVQ2SxPS8XKRIE7f/ENrY+1sPxVhCq+sgVYvG03aXZJQ8Wq7FGRKBb2htzp
4pS9Kk4ZCSvVOtsTyRBT2fSHqtc9Je5C0EB/9zR1hMqsAXj3o1WaqE0f90ntC7kK
SGHKgoWoekq1iJOvPCQvxAH9JgWIssejWATHi2ViCbXJyFQkLT6SM9wRgI5lRAYn
LeaUqrIK+bYm3su1iM21t9tTYcPGiCuLtq62U/HexQIQeFddkTKWibHfIiYTLtsN
d3RpsPu82e5OahG/V+kT/mzKEv5+Ci7DHPXPCR1wclyYuokF0UDwnLn4+sUTF+fQ
PEacJSZMmEbXbzsNlnIh6ivVDi+FBYf2nbqLC15FCSR9b25p4bZV+fcV0e3A1MUl
YyLYnJ9oasDTH1d/4TYgPm+Z74eceuo/g+lyvCPudFZLYClP31FMTnypZbieQcsx
au2ao6UPoHmP5ZCs74nlJbEzAMMx7a4iM9vcCiLIzx31OqqfYxReroUwb1Mrp1Zw
udFg1wcCi9wuL0GeJaivmMilwm0+Eqp5kNfjDBuFYbesO4BDNlxHfxqFImpCrIA7
p9gVGY7+n80yTCM07aGJlwQWk7FTs/JBVVTaxxNe6vh3dsxcHOy8BapQ3ZDd5i/D
kdOsAQu6z05sifwJNuawBSczekFM7BxsK00+O98LGsAcQK4IkqIaKHq97RnXtAiT
gHzCId5oHuUso2DHnTY99PUGb6RP1QEYLRqPMFOmtfaTG82K/wKd9MtIOVD7oXbV
DjfDTDqvK+d/wbGOjiNHzyGQWOoYd7dNYvPdlAX1Qh6o6w2vqZwkWlyWCfeaEtSB
L7475gaqU75vZjvCPZ4lAsZVrtYDCcn1lf9DkletlRy6rRyfmP4qq6012zhCYu4k
vwZS/wIM4z/1XT7yJqW4xJfIO+xSND3nDDN+6JfsN8lIZZ8KLaXoteph5+a8nlJf
j12Tv9THjc7li53zW5f61xAkUVdHsP/4/8WHAols6YBBsbfJIRtNtacKPUQyh8XR
LsPYAmwMOoYRysxMhkGr1/i5awfV9mfjOUem2aIaPDL4UGUd2xxmdI+0ZqC6IbAx
7pFTpjtL3mgBNFXh8AhFQT7Pchl/csZdZOqlBtqB+8qg6LRqKxia543zm3zbQKoY
XVrCF6DwmAfWS5k+ezd4cBkNKbYzSV4tBNiyCUpg0MG7jkUuJ54FruAHl+547ZjZ
WRcmlx1txQ9Sl++hz/a0JJWaBho1f0OvX/G86C+yG6xNt+m4CmQWtjhVbCJU/uKw
03SyjQMJzPLg+fzaSPFH4bkhytvk5f7RVP5TKCgl36Gi0XlEs1XqDPQYr0AePD0s
5O/EVxSo8v5TWydeaufP79JfPlmWBLBpixYTOGoajdf/v8PQDfr0tRp2RWA7BtaW
snTOq0iGmU+qbChqVUsRy3m2fE32VXDEaXmEzG4vLoqgQyTEX5UFhdQkKKPEzCjo
oDdHL91exkfSL3oBehoe0+tBqpg/huDZaCqvJPQEBE1HhFtJVuKWo59H+QamONtT
h0zTYTrCHBw2JbysXGADV+UveLyJoBeGspJ7Cbeq1LafHrx1JxsJ0+y7IVFr/Yzp
c8P39UB0ZsK9R3Z5aq+zJ/ebIagSSf0bG7WP+q7MYusoIR3wlKn/EoXK3bk088nE
TmQl/tSGZVqQeG/gRF1IjKa5yCgiAcFyJUM9VyC3BgLmZV0IEOJHPjS4oYmNpj5n
zvoKfPfTsou/Prv9OX5Bdw1ZWbxe4kqZqC5g72A8D1wqzJ8eDlmL+XGJ1fcOUS5K
/HghpfQbhpdjLBd/U/m3QGJDwKGCJbNdXD+mxsAv50Z+jvGmE0Z8YNAKzmj67V+u
woFsj6BJ/7juTCbkSQ+heVm/7EOyt9a0/MZHoKZb2O7/sukZpODhEyTp5Skk4qPo
xJmqBzJ9DbxLZHa34SrdfChcpAhYN0jCwQxGGIvGqoFXDsOX2CEW4WBHSUWhFJxG
QMkV7o0XYrBQYuqUMrePPoGx8GZr3lEQ8+TPlt9OqkyT0Z64jSlukQRD1Ufb3Yn1
msz2L0atR3+7S8/iqwJwJSxjsosXGsSAm/3kDblM/5J+9cRj85e28wiE2xWCUNHn
lA1kGG4Pmzj2eDkg8NLJMDrT83dAiFFCF+p5vokSBLBP6XQFadUz+rLoOSuzWlHS
UCeOw3croKJQRc5Q3jCe4Wg6PhpFs7kJ9p6e2nsWcYL/LSS4H1wW72YaYnp8sIlf
7meAWR/dXIY0nf3EJ0bs+n4TmL470Wjqef53/kB/xwoYMHdkXmm9IAV7RWIoTREh
UDZQYlWP0WgBQZGSsfvuVfU5DGiZdxSv2syeDGDu4/dp0hm5N84Y0mkM342PpRoQ
yahANC5aVbT4+a79zgywDYsjYpXeiKQrbVAJvXkkxDaV0r8YcPdYWVhvleBMWggU
nY7Vmp30AsGr2ZzyMUlDuPg3qAdR+jVckqihMeZdFERdRqpOfyH2nB2kM2Qgzkc4
XrQiJCNQBpygNvamXolclzirDax4X3sdjlqADAqKwKxZL55TKomF7snNQ5xF6ZIl
DmoAT95D5AXVySq7i/x4Az1SlenUKjKrD3pjzExOede7CMrFeY2fcYa+Xvgiiqi4
F/vxEgm6MtS4fQZ/qs/tL2bVKtSjDasXFlYBLMVOmXlNs8IyUN1ibwPMehVe94iJ
4tsNrtyT5MwDovz7xPNW4k/Oo7oWomUwVQAhQzNdhDyGgA0DH16ofNG+lptBizWh
lx1BQiZklKb7mzsWyIMt1IwTFMckFv/njSP1R2sP1phZLjILsPV+ueGLAwO9eqtB
YR5jtyXfb0AfJM8mFgNE6EMpQhLbXH7TdKlPHar1mZcpeNWopWtJrGxwzsYTdhZF
ySrbEeK62Pb5TfzvYxjiGEDeq3eqp3ek1OKjip2HI2aReMsezyXs4wDpXMaKPUUJ
FP620KMqLjqNHEGJpeupwndPCMhYNcDuE/e5TjdoN5DjaXnCtPl/oqaGtKZk+8//
7bNLjgcMvMXZH+UapmYlnehiWG2Iy9hWQ8jkfs/A7/FJCD+JCIRBt+smN4l+CyyU
tlmNtMbI/nFVJijO5qhOTKek7Vj1knOLFWcSdrSRbqRF7jP3ceZeebUmwgJkXz1u
uhmX+nd/PNT06h6JwXhy6uPQ7nW2y5kGAMVU1Kb85c/PXnYy0nr2QfFA4wXfi1Lu
jg5O+SimFCRewjilvbOOvA8uOby58PQax5jE44WhSL4Xy8Obmx9JdGnrhwfyFip1
4P814Tm2hU+wRy3mq9qpv+h16zjG4f+8eIcUFyzqcscAinmLrMvC1IYGoWj2nRSB
ns/vpRp69SkU8gDByo6txLC98Fbj7RsptRuj8NwdzO1JT1Lvpg4wym9UuU9iWxYW
//VDD+r2FBceZQ1PO7ADrpi/OZZLge91CKHLshTLDsZeTrAT73FBRKBTBe/wDzYm
h9JouVSGF6ldo72fk5zsWbgJMUqbZ7jgTv0KSfZYiFOEkYyE+Cv3TbiFkqXExTqv
gob5H2bxoEQ4hLQgVbtj+FNfDCMlKcX8QebpVCVU8lxcMDUCdJ7NzUc6/XIg98TD
eHjpzXfW0SfWH3jT5m1oq0/7fBRUb+at1Fl/dA7vOI+teYXxMNPfP0jM63JJ2gbi
oIGg1rVSlW25y0EyiOo4rUsGLJ3Uy7t9X2P/ZGS4ZTqfZoIk3w/TzbBdcmPmHGfh
7IoNSd7c0qS+6kv9Lc/oaS+2U/CIGifZOFAk/W9vcxGN4zcZggi0XNDdgCTDqrZW
NGJmau2v97GrkerwUGWcIXMcriBdhz2Eyjtk0V9n/8d/KAy+TZ0IomyuWeeaz7yU
/w/8f/5Occb+3cO5Qt9mq7p5WS0unCCCOdm1kVmfxOgmhxDZ+XdRRZxXs4dluhWm
TY8bqAl+BoZ2YLxq2psM2D8cHRnZU/x91dFpReccLClH2TNP7Foftukj3zxpeRzL
Qy9KOXvo3AzRkjr1yBZP2apGr+CJoFhF3RbjuKtfGI9Fk9LVGHuXqzJgKCQrBhPY
Waya71cRydBxUDigr83U4GfuhPJBbPMmDrdQvoUDz+NNrdIjK0at1OwnzrhG1dor
1+9rb6n+/gBjyMeMeFRWLu/SsiU98dPecYtZJlqtLCtjhy6e3drxpJIjQ8F76xCN
VSjsJuia2Foz5d9wbt5e2wpL0rB1nFRyUuL5CHqsEstmxZqc4iarEUW+pzUNERq5
2K1h4D/O5HK4bnNNDFVfKNlXTdeleJyXRRo+0jYtRXEi2/D/X4hen29/hxSpBcgU
su2EF2DuITl3xlHjukE44ZGHqWQYRUgG0+HXzsdlioZz6ZYPNcZVkeAkfqy1zAlL
K0ymR3gGr9I4SSnN+hcmBCtD3+OL7w8VUadaDlG+vOD08xmxrFB46Z3u/6th50ew
WJI2D17H2ftsayXbPbN1rzVdectWu76kphieVTgqpK9SfGu7WDe6artypUdhJwZ3
hB4Jw5llwwqwN/f9glgQcWc4ZQdhgu7gX+e1XWAkqmuY1TZwsY2BHePOOgIM8L4c
DVbh35rz6nG3sbm53nA2uD88oEhyoxhz74q3vcZ7z4XDHmHmEv898vIFpQafDR24
vcK0jpvQH3MQwVhMi3K6QnTaQ2lS2/Q/SSp/5jL1Y9l94F944TMWZQx4u7qEaZFj
MFv0RlHAsJncPXKCkntSxLbgMswBeEZ6DuI1bTn8JLj6meM9Mu6L2qrbmtQ5bH3j
vpQ5r3uLjZaKL2+P/0peWWsH8aJtJrs3IvvbIJtLUJ4p79J/EQc5IwAvgYuOboiw
nKvlylNBjOp0ivQuDh5N8DQSha09eKIaiKfa2T6J8yYlXgBf8DoaARSL414yB7X5
3rSRMWNgsmfV1mcGXkOsnwhrVurbkySco/gKPRaI7cIWzXLdiLtttFgsVQsgJAWN
WsW0/1uNktu6w9SEYEAcZB5e0p0ZXJQJiglmAb72H/KC2QviBAoIbHnYfRHFFkWn
ej+zL8f6tHN8gn28hTrhy+ixYjQ+BTD7BzokUZxRO37ray3D6H18PSsRw8rqDtYd
rpX7jkpsqst38pmGE8kf5Eh5Pr9AHGFWkwA4TINoxOg0WwcJ+51XQEsq7eRltiFA
xSmctf32pY44GpNrwY5ouKHJZey6B2NL69XuWm1zQ3ApU7rUMcjd70OLVUA1dXYq
eB4l9WRg7N1gs+RfLsYqHuO5XEfmrByQjE/GvtaAygJ9XxcU5+x0OC/oarlvOm8E
HE3qHMHj1qETX+QHqLYI+w+aq5aI45ArAlNJ8agLkytJmzSHuVNRQDHM6ZQq/PAa
eW6Shani8Mv5n9OLtQigqYK1GGIPjx4Ok/dAKPh4RHzdWBzFJ7CuqAEdvXBdI9yl
ThCEkv/SOD1yeHm1XU4eIyNyLG+tglFImYKRV+0RZmAXQGVUq7x5NFhdYpdmMI0C
lLnhfi8bSdm3BX0JvWS/gE+/zOhO5DeiqerA1cky0rcOi/h+E2CHqEZn47hTE2iy
xV2CQyEI3x7L20unt5lU+6NkljYDs1uA4BX+dq/NJ5DE/ydOlJjP3y0t0f+nY7ag
dwBSY2yr2TcK4wJhpeHwkj6gkgkJUhKUuRMXSFjrZx7KSdpayQAAuf75CPps1TK5
b55c4qBc9ypOEBfx6PvI7ek+zc1m9Xql7luwJt1fEHSM3kmuODOISU/6jgcY1lJw
2DbPgnWRskc2rDPsxziijaiO/nIKnthHjOgMPvTRx63W+Cdj/XNKRPc+BMVabkY9
EjboAu/U+Z2967uBRgQW5WCHVH3W99nXQHfEo/VB96Xf82qnyprwdm6fZhb89s5M
a5y/nH6ACnSJyM1eKdiuc+j+DbeyeXSDKa2GxzcODv2JwA1zPBYkF4FIsdV4qFKc
lomal05BdK8lW800pBrujeCq0bY5KmbSSKmh0j3MBeKLqizyMWFD7l6oXJPJL+C0
lSZ3vGhrMkfW0ehSTVhL3WMkhsQjPcYdsf6HmPyiGUlWr9YzsCjTLlD1dVepLdeO
qLN1RqHb/VWyQyxYkxyzG7XvpA/8eTcBncefxPCrbZ1a0ukQb6GOL9pFjMz66Jsv
LJjvRa/VCQBB+EVHzZWRGA1NM3xcpQZwpcyinzu8E7654FvD/xVim1XOIp4iKlun
hYDyNCkkLy/uCcgq9TBMUdAfijb1asHoSA14d2bBlHpIYP0rYgJ6UQa9OkobdXWd
LCha8Ou9z5+pDhl+PbzyGv1RtRdB6d/KRuZPcnHzpGHiP4r5RaG97m1F6b4Nw7nA
v+QCj+wqEZWhJqbprget0mKWwDnXwmzv3UaNQBjllUa9UufETdyVADddmuHSm93G
xNAP1c7jojwkHg9j9eXjqxYNkA4rZ3ZDGUZbw/GW3poAU/nUaBSur10kvSj/qBHN
hh/FaJ/JVkWNr9OWk5Liqhe4utsV78kRjXuclnJudLKfVeDFQk42l/RCDQyeQAQu
iG6HPEsXQuO6kvwG1PTgbnc3eXkrFJjxassaJYFTX99I238oEXdE6etRkzYsORxC
WO7OX0n5b/q+oaxhJMoDW8PlwTDRhCPdf2IsOVj0+OnVvIc4mVosF5rnQabd5Yd7
RJBDUCowfjAiqtF0ycMe8H+REKqfepcm3sBsskFhVy5zmVyXmMc7nbX8LoVZjKmU
t4SL7xuaKMDTpUAfeMnAS19pqdJzHhxaUWOMGj7RKoZIqTRb+OLnvaqwmWTDVeQP
Bt8WbWT0gHpprb48+Zf1Pte9vHX2Vi5tR4kakSLxDzOGVZlswK8WsRHmPWArrZPS
V7jsZxL+o1+2eDVCEMSUpJeiHk5Xvcv1oioUgNVD7Wh8ukz5hWdKKBQHaQWo7OkV
Cmub0wVH4bUIAcoLN500qy9ekonURaGRsq2lZlJsen582Sa+dEMPvP0abMPlk6v0
Db6VHzHoZlepga9ClLyvuIIfkXll4a374QpqgfPcZfHLVt0PyJ7MqBgVrhpnWC7q
71AlWArjR0/x4inV3qB7lh4T+beDt6VGOEKr5VvGwgDXUlXTDGVf7Sd6YdKXXyN6
K45wD+Sksg5VCHOqA0qxEAJ+KG3uX3/56B3IZMWsDsCDMI6QmHE2bjW1NO+ObjJq
YjXzuZIi42p5yoxMJUGLP1p5Ms+HCO/WuYFSxCNlrPNPVyQFLeyP2L2pZrRoMjl3
L7m2DMDg1MId2zNiI1DMSjr4Gw6C+wZeu9bEHsmu6c8groewDndzJvG9BH3eD4Aa
LgiRR9LRiQadqi6do+APxhiuphyNyNj/tW5NVHtXfsiqRkgbNOJr9sotHkvOz/pJ
iaPCMQ440zgfeJN+art5JfwP4JXTUOVHe1h392za4Fp3LF2LwANPsCDVxiKkdZ3k
VqhNRj7A1ocSRr5cnvYhzWbPP1fyRzASL4fo5w44Qu8Cgou7lCnhmtwXsqzn4b4J
6yVrvu1wnrcmzcpyPodjwE3qOSBOuHbj02PBwjOpmVD+2S8c+M+ccwKtHUY1ADIY
6cTpGfftukdwD2eFrYDiwNoBOxBA3gIYm1ywuJLOCpsqpdvZGyJqMPRXtXtmKEoW
xhauY1tUThnH/rmeZUGAygsiVMbKQBd1MmSFbtDdsg5N667wZo6iOQ4GEs1UwCVQ
l+uk2vuuTkctesuiuOTvsdQVLMCZ/g4FD5Rx0DRBPFuFeshi3o1vg+SPzOVc8AuY
XZ1Sq4/V65BidCNQ1kCHDsUBEph4c1dm/+ySFfWiW46zSWsPgG+zGewtBN35TkDY
fO1R58OU4ch3i1TLZooe9/FtR6xCTqCYMAjR6iHfCjs8bJSLitH0ji+eptAJKsNM
c81/h5g4Iz7eZc37nRtL4fTLAE2iTJGt4/mX9Pb2UPTCKPNM5dq3lomMMnOBWc+M
e7WqKvPkmFBL5oURWbXsVN/dSYpExHP9hYXoAUWVStFOP4FITi9TJ3M+O8GALz78
cEQ7c9Ydoql/HUHZfT9qfjtoC634up/mOb+07HhlqaNNHgKcRyEuTJshcuE7WLoX
kFGzCAuaHV3yp00Zr3aLpqajMsvdBeyEmuZh+y3r3D816rChGGPMQoJYb832AxYJ
b0QYT4jTuIlzq1NyDvuVlim6oJFOw225E5bT+J22lDStUEqgiOFkm+so4Bkzhxli
v4G5XBpeTLr74PvCRqsWZKsuk7SwJAVHKlRcI52fp+VGT0Y3SrYZxoZw4rwiHtry
TSU94VnTH6rCxgeUoMK5cDLBEigtOuQ9hc+ai1S4siMhtFTgxKIWd5rx/U+Nf6V+
Wrbt/Firz9lZfenIeERtCUslVV/nE3jzehyqjRAwGfVZmE+XHY1CoMUzqM8EbKII
i5jILyfjqyzhFlwEGVnE4ZZwSE8ik8nT5qw5CJSUcYvINJR7IHY/+Etv93Gr6Gce
/owWy3uvhSUl4NUD1IHQnv5RcuFeBEreVe/Ty5ztY9cBr5BiMh9ZgBz/b1WU7ptM
//P3n+bEHHxkVWIUB7GjVc5ZNDCEO5HOmrLl6eIeIOo5aF7aeig/LA+wB6t6sC/W
5hV35wuhVovAtfANxb0TiiSrFdKM/NWoDAintrxKK/nAw9mAgL52njr3ktrfrhkQ
qwvuc1rGubrv2VWZJobGRi5L25V+FOv/zrshSTVR0pba5Pv1jKi0uBHTK/l3/DyG
wiwkkByStA/lmLBVraEB+otuupR+yYolaAdMiHJ+jHQ+I/PyoJbdTmLuUWr8aghF
8q+F/l94V2JurqwJCXjX9DvTCY2Im+uOOQePMI6D72Ai0a04YE6xvP+9sVGmHV0F
tDW4husuvNqevhco0qJ1ljVPSWOthnfS5KZ9/8w2bY+iQAAjyP6nRMWss0ByzXuK
askjKBjB65JkeC4IpV7APm6s0DtsyVKruu6CBNkm9ov1psqPfc6cASBY+dIuiPHj
4GF0mlh88yftq1+kGe9MCBI18SW5RcvSVrlFTaGT53tLm3fP72WwToJ0eLBgGz2/
W5tgzmZfIl9TFXhP2ObEvsQtPQpqINbOSPoH/VtbCmMF2JSIyRWD4cKEZV3h9oxe
yQTZuexmCPIeh/vcqIBox9UuXF68Bb0Vdrn28EIJH8sRYE5+yiLQ0UKHokhyfyav
D1Ue4YB2yG61RHvcTUcDEZI4n+1eF6wR2LSZOjepeb9mIQhCW08IXcC1R1SVE+1p
ssMYMi/Qq8Mh+0lllcvwzA+lp9zUzuOfvruxtVvKi0N9n+0/0pm8/YHqTJWz5BnI
XBXWXDuaFfZDLRAOfxK4fIDM1N8i0QUR+xsrN7oxtX6Q6uki/ZpAiT79c0dz8OEa
foG+uAgIi4lveqk1sCiKw2OZEqtr+Lxrk2rBxcsq4pDMa0bFO8oQdQfsDVqn0LNW
DozjoXrptuUT+/58jv+CIiyBbiKnPC/f68k5cFkSl89EFVastUDXgLLrdY9JUI4U
nIvssCZ4xQsiH/6d8C/fhvMrZcyLT3TbzUspJxGHiatUC4ln3UiHouQU0ZtD+NfS
3QEvmFVvcEpIyN8S2ABQkzgfvBxZEHlxkQDAUC42DnGh23yKiuuG1lv+5OsXJquY
tv8ok1pJFzDjJrsW2+cn9WRNIi9kdiDcRQwa5qA20MeeJxBeCq41v7LU3ScmkAdm
2QAxl49n/IXmiIoAIqhO30stj9jJfNee83kPDRX7qZUfn7MPSidJIEJ9EvaQoe77
pTtHsEFBu4A+mShgU9Si5L+E4wyLFeXYUjZeDYjk7N/xEWxBzFMuKWQ3lvHCd1Kw
dVihTDsJRnl5af80BRgp7sg410TzZSJtQYK1/mSQeOCCgFHRJUj4/vS7aM+OQ9Al
0bE1/Y2aILeiGf1P2gCaP5dYogYznqbOJHkwBtys2g0SMD+ZQQO1x82LcbxJnSW/
CFO6Ez0QPTwcNeaWcL/ngk3Ia2b80vqpyvH/Kbcid2i4kMdF4FNBd1T5in/V0Uvm
de8C8fniL+y8ATO4M8+Vjc3l+8k+4Yd+r/DKbrt1VIIkNAJ8azgz58TTtDgjhwLO
T7fhruQkmYm3IFUj2nqLh/FdKTVhmH6Gc7rDZUyBi4h0uKx0a3YLxhsam+Gl9b36
KRB3kaVGaPGAVgQT/dpjeA/O+gskNVI2hdbmz5gjefbggGlFuQrQwV9r9XADCwfB
GLChTQMIkKWuypn1jtdhxhJXpX1whIJ1X5Phi7I3KaW6giNwlSJ67LliWmbYTV+d
mayyBm09uG/yDehshrgY9smwkuWl1LMp2UuA3RcHGBw4T1eKzaLES85v3BwzBnaV
iZUGpZoqtePEKdsLJvwqjWIjBSe6+AIlW1uPg8JTKOStgtDymG3nrm58pA112IDS
PLbFqjXb49d+O1Az2mS1XIXwQ0D1t0I2Mr6UnK8tAd30/VLcAOOQjMGQsmYKx5HR
hy7e+kn1WU8qbzoSsd2g2tfBUlGFY1qj11zW7H3aEmIxH74U0N6q8ZsD+VWOundO
Vs+/ggO9eWFsqfZ/heQRyPbT9/rcSY803fK6E8/pWOR1r8fKbmc1ldr4HmAug3J/
l0hIYJEUrh4zrITBdnzBe2snSQFzre+Bem2nwCJUROkqZFMuN5qtL0uz8kcnn4al
YPfQk7kx2oxya/pl2WIfpHXVfeCl1qQH1VDu7XnaXLDYVmojUHEq2Gf9xjTIkgJB
yR1JDMZhzFyiIRuC/I8jg2XTpP1pbJECIZAx7aIJG6sd4qHwvQK7myDGPWxb+O90
bBuw8biQDJjAX+Y/7TFlGuicwUhsoRLiJmGbJigV+rajBWkaVmLZMXoWB/CgPHMb
4Ue8Jb8aOf9ceaLxkGxdmg5zaPaBWxj72zPOwUhnICiAeyZYVIanEis6rA2c5Rew
GAYwqstB9BUkvDZuoot7C6mbPtrHUBOtMcuoJFhI9Bi1Jdzq0JGUCewNMoBPtibD
N2vHU41tlF66dc7PGILIBYuyOXIhpnxcRcnNK9IF5e8JEJxToNJXFBUpMoqJkBE1
xamT0AFu7zX4cu6ixfuWbQTdQiXyv5HTcP/+3riUi8lJZ7ugaj3wiZpi/WX1aCkw
34Hjsvxe42qKEtFWpgCyMP/hGA9lyWZitzI1wCCp0RF1fbEbhvQOZlWr4jveXtN8
DTAEyZhhnkLsvT70h+23ay3DTd8vm7CxLumPE1/V1WI/bJmSsx1E0/vikAxUWjZT
KateC9d29sj+3h4oF1reh6XXSGo4AYiu7H1MQbNOSQSqil9bTwelHww6cI3WIz+H
6mmLYylvebkNGstdQlB1oP2DwpnqDqeHnOEfZs5nNcZ8ZxOwdAzIFKrZzYnZwvGT
zb28iDw9DO5dCVys14dQnZHMtGoXElVCtgDaOaMOTnvZR2Qjlc+wPFYdgP5zB5CR
bKnOY3lOu8ptHv/nqGr8l5aUCg4dXVbTwfj5xFIcQMm4X4j4P/byf5dDQZeBPZQ8
7i7M+jQ9c4O0szi3eas3HdzWzTQNM2v1iX2SMMnb9PIoOVWMm+BVMNB58XlpVs7Y
5y058NG/WfApY5vazR2T3Z5NCcwbdcl77b1ZPIXhRhICk6Jd6mK2J83oxCF2GPyj
y2vUtb0ou/vpACorzgukldlArXfSn4OiyYgc4KYk4x2XVxZRJGK/J9AKTOGfS0xy
DI/irFLTyrsI4MS78tmFG3gwvjaNJW+Dm1uD4uPoLsstD26aEJEmis8oQdPwJYvT
vaXz9JcVGGyzMvturWi51e3CtHhIUkSQZiyqzdQv5LOzSenpeA0h0IjjeWNtMp7N
KuI719EAm/Jrsp8r0IBue5Hh2PydKxqL3PcyvPARHQd9Na4RRTVYzBOG1KffUDwx
yNEPi5mPnulims4F0OUTJvuBL57xqzwJSgjAtrtjXUEBMHX+vrrk9pS/VU2BL7Pe
aet13Uo3wkwY0qRYILaKxKQBpB2JHXFj18nIYMdRA8tITT/+6roTPjVi/DLL1x3H
JI2e//GGCAo4g7isXQOPItiF1Q4YSIQYKCKpTgS3eYOgBIPOmtVhYbdxyrxNjfXv
Ap/zUIshREfzKhtFbwKBUyB5SSiKTaUAPbCdefGD+X5WwzICK0DjNQNFdcXoq7CE
ziM0iOlMsHQlO5F2OCm9cey4YBIzYcAGeSq376oWyhzlp1BWy6MCfGUW0hgl1D7C
mNwkxmJrx80YlaQIcXs8ollZ0Lyhj7FBGDpUWpbC81G35wxV/Qzs63Oz3IOm09UG
zK8gBk29aFJaR3/fv21dbWiDfvnY2f38CKQf5IWuvtqXGjKOcm3DqYX59RJ2A9fX
T+4lXI4CIPTBlP9WTGUMd4Anc98I3c8TwmYqZeoloMVGf1V5kF5izIbsxwxt12Op
QjpGk/f7TFhgzSKc1XGfUYGFhtA0m1bGMj79vq4Qknhs7+a4tmO2dZN69CuzOVfp
179jvCyVPmP0IZ6CIi0bCe3UFLxAba2axYlCm/sdaOI/DpnAfMXc8AklK6E60Q0r
ueJ1h6IQl463KKCaro6cs1B2fkjRHHENqo++dYzp77GcKxV+tfHFrWKDubP3O8Yr
0IPSOCYVsTs2z3hi+3yaR1BzKKTJHyVetrVPC3for+N2JS1hyzbKyPzrkzrw/QG/
Moe+6kA8mk+Tk6gZ0+55ETIYnzVAxvgr5zdqrYykDSmLET5WttxKzpyF5gtT4NE7
fqHhkUbboZ73ApuY6rmVgD5x2FBWhZluDnEjcqg25AWf1QqKRgDIxwfj4vVG5+9n
+o+Ti40LjjXp2DnqZCfFDKZ/KFGU8l08e5sZVfseuYwckDgSHifeRn9jw/8L+9EI
uNYz6vZ3ixW+uZ7UhfhQk/LSObPFVqRXl+jDmwXhsrz+gngnjkgNL5iVija+d5yh
OTlv08N0mTla/7rg838ARtfcHohW7jGF1wWUTqWZ52uY/vkCRWLmcc5Wc/5nRWI5
nr3W41oJkthwP4FR32Xin+cSFDwGjuuZfInGi4cdInXTd/w55W9YLEG/v0UOk2w8
bbG5VrjCMyD8XxPhMfNOcaEVCvkDXkarPALt37K79HkTUWvqGgeD7R+2s8REcKsX
UYUAL0S2OPdIy3tE+FKbm4w+09jDrAXRaB7cXGWhK5aIFL/sMi0G9PzjI4G0Mokj
74IoNqXK/tEsqwlTEQmxbsh/VNajRwXB8nQ0+t+mtIOkuO7bdDufFq/RXNh2bi1U
+Sz8vpWK7y6ROm4XS7jGXMhB/u6+YJAPRIxUhD/lNtWZanDTgKolJRSkuZUQVPeN
B44VzLhHm3Tus+FvVKtWsLcXorQyfmGtDMPQ6HHLc21xmpXJT1PjqI7GIanB8ErJ
gyw9RPnHyv0CUq3wkmE7XTJcLB3xdMYK0uazP4548phDvO5h/f7ZycpqjnuumGkZ
z8c40Ouuo33lAUrtAgTv8CsszJaXJdwriv0QIPyX6fSERAuJmHvG7iAktTZiToBu
pIvOUZwz2DOhdk5eCCzxwhg9JIWh0HMA4RhkptLtS2serlDBX2GrMW1aJUh+rHQZ
IUTtFQ8PLTCbMpzr3qu1MkvoTOdfYNf0FoIFFaKUNlOMqma3uS4s9aE374YpEhdX
NPPqdMq7jhHasGiuQejE56ErwDoZhPPgmdpdKmaM6LMQfbsquwUUm6kapSE3xq9w
c0rsIxSmBrs+xjphuaRJ3ZJmH+FZ2CKPQHBG6NGO4I7/n3/YX9lYpNK3OqKS9BQ7
IRXu8fMeY8HjRbj9Bmm1uLjLDVdqGz+qzS5id5qpuscDJXQwcUiSwrV1rVxNQCsh
WdmlYmsaQzi+OmmAPtyRBr0hKuwhSEDGRKp/1eRmH+3gpWzhIUTsY82zJHs5aUCo
GYxTsOLwFL2gA4AfudpxflG39DIBjqydnIhzqzT5xtQtMQW2h7/XW8A18oWMynOM
SZsCB4zVmAHcZ9KoiPJl8AP6RVrXgy8sEzLgkuuZ76qv97RsrOhxn9kv6TMKP0vK
4wNtfaxYXfKwIk9kOCtbcI/Bt36QsR7Ac9KXjo3CA1h1N2x2GAPAv+gh9qG3PT0b
i3Jsj6lCKoBoiZYp0mT19cYro824bNncAa9if6J1PtQV+9ZoE8DqiXBRDl4EbneQ
tRMkA71f8wqZDD+nCqn/77aK8iXQ3Vr7ioJPxu4mDoxAKygpdggdVM/qB6XZoouE
y54Fd/jzOxKgssdpwB52zHne29cIRkPtXaMkOb9ecWHXYVj3LoOKEIaMnd+y1aim
KN7qvDUfmiPfmojQp++k3uh4IQyYLN2s22oGKWbwP6LDUz8+kwcrDYfkShi0ELDF
N5+OE9qfHDMfKepXSuEHB2saU+z9NAyZgcxI7Wqg+aQRtDWqI8ylM290z1j1cljj
NunObzf04M8PvMlK/b6Ibr3eC0d8wSfIYU0XCJjvnNnok777mKyAgFyFBmkyCnUv
t64KVcgP7gPOGk3uw5rDtgfIi8jpDhOcOxIuHogyyHVSvIia24szhZci2hI+umUS
bAgL0V7EXtzlcq4uAIwxWlCiCI65YZ3qkVe6sQqkVk+u8MxNgIdVkVn7z2dv27dF
pFCSecbpicHivaEekMgJK/lqnlNiGKCpsah2m1O6bzFPhWKhF0k6nUtC2eT3OrPw
sZNKk2c0NufmewXTs+VRleARsLnltXlk+AszDB504a9Gx0Ig1Lh7AvEzyspUiTLp
R9o5yu3S2ugjjgsOXSMy8at0x4sxzavdnT2J3dtqgRi5SthGf1vfdPCMG1OJyB+e
s5kOBAnS5tnvCDEiEFwscqUagZMFVwY3Z3w9+KAZyya+1Z0ymeehZcI36ZedQYQ5
6OGJ8/go1GnyMNdwkOfo9QxNGSp+oBwJHqp5dBFt77GttUuc9RwkC9tqmqNo75vD
oI21m/JA0AXt/D5BAhMTQ+noJsaibMezQOHys8rf/X6Fni0ocAnA60xybUxiEPQ/
XA6KNyDoWgSRKEmpxejZvYkPtb0AJOYknVIaGNKpw/O04DtU9UsXumk+ORnE1k65
uHhfx5G8/ol6Ihu6BlCAhk44OPAIqxbGmDRK9HHmEx1s4spN2H/+OOQyFlNrCaNS
tuWoDbyrzsB5CbYNtCmbvJcDSpqYaOR5sOCLKBuk2cYKpafWEDOdZs7r4yU/gbI5
0Jyw8bs4XrzKIEU0xVq6gGPP+BBDlxMJyyvckZ17wSjDxe0R+/fHumHCd84URHWY
mebfwh4fojelaoP7t/UH0R/24XgmdnfjF40BQqzDUXzVwveeyCvb0zB9scEMWV3E
SAvb2UD+iw1+rXsorSexHxvhfArCbLuZrq+Sp6agD25rdhuX5N9Lkb6BaXV93VOL
o9UPOh2PZOR4SZbkFQG4wwmV/e/BqnFt1bxxwswc3Tw7Oh9gLXZaSo0pKyz9SGb2
VD26oI7jj/fCBmY1E/Ld+9Jrur6LIpoKpLo6xUi3KirRVC5PlMyLWex9l0I9UoOT
Ws1pYmfOc+3BF9/RdUenApI0TcAVtFWgRNvM6H5lV8G+UzRHi/LEv8tjLD9ALC7d
xnanf5i+V9wfE5PN4qwXjjmsTcsbbR09VxSJN+fSI8YIjuLeAKLbkjwsUrrKDKjy
sKtBRoHHLEiitWcPZT6uYhNvGv4V7s0zcwzKESf0big=
`pragma protect end_protected
