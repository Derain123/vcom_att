`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="galaxsim"
`pragma protect encrypt_agent_info="https://www.x-epic.com"
`pragma protect key_keyowner="x-epic"
`pragma protect key_keyname="rsa-key1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
KaTG5bUH1J10Jisy8E+TDH4SMkW6tESVOzeBV2OAg0mtVJKVmCeeF/S2j1W68dng
k0GRVGH6Bn2ZJWiOrE7wJhMjq8DAccsugbbzTC/t0CpbPxtNqenGz3j8V0tRQCBF
75+vPwiuB745cFTqGbRY7YvVqUB3ZZVjuZe7aFonr8wb+2XS7DNuBmInUQvky6nU
CpPpjBeC88u0TDGTDSSWF47s9pTCoQO7FKc4b+wpor2ZCA8eUqjkrulbRYcqtzM9
ZtwZIDZwJ5Q9N76Vok4qCY1YGbl3evOHJ4+TsXmjrEKhEFhmVGYu2kWksTlaxHkA
j1PjEhaL/jvRtJQOpdi4Ag==
`pragma protect key_keyowner="Xilinx"
`pragma protect key_keyname="xilinxt_2019_02"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
Dp2n8p3CmsiYplpIGcwhs0eXXGY6AC6h1/uXfmRP+n6d92QUs/eAhpQBCmVdbub5
4LEEj4oPyBB/rQeMTdiwejLUskxV4DIe5W6SSrKd2c2cQsl2lAOAeWinqSENIhcl
aO22PK0LzFIaAYIZlB5Z2X0YI1QCnkIJo5kx6ci9UafyTdfnNaDdH+FPRROIQRf4
tLFvGLOeoaW1Mh2cQ7pMq4j5xmkguWSZiyJr34mSbz5r89Hf97QPwvTEIRVD1tvP
tmTIpVX8lvfwG5MZ+igs5F3756KQEDuOMAyytsispU7qudrqqYEsSPvasLkRwLEi
uOq5kYx2AlR6w1Wagqy2/Q==
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`pragma protect key_block
t/OdwHhr5SPQcTeGtDKAEM9Ml++aBjlHZ6Khywc8InlUon3nV9lkFt0FN/aWc3LG
ItSKe5JUoh0gmNjx5sYaCfNkYbm/Krr8vSUeEoIQ4lBLDxf6nHAW9X3lVwaKYPb0
sCvJP80oRe2qOZfsyqv861SnsmXPI8eRZIW+vCvcnds=
`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
Ub0P7+05YV9YJS40hcXUj0hni06b/Ur0WHXw0I6WjdrUL019OkkUJlo21ohlCNFT
P9KnzL4XmXo4jzI0Ab97uOkYvOM2KcaR+XWDMFlyY3QgqP7dq/IULgpAmHZ4ZUjk
6xKk8J5RLE/6oip07OrxXtOSpbSaP8Pa18xBfQFmZxkmq2Ge4XGtgDP9gCbWXTAg
5e9Q7xKDKIfZzModYa+LOdiGypyQtznRnGnGavSPql3+v8nsEt1keObge/zfMszS
Iq0xYTPHyPnBel1N67fRXNghSR+KkrL+9mz0Q7Of5ysS0FAyXX3eCtx9WqoA+UFV
DFvIR5Lz62LquysJOpPJFA==
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP15_1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
qdSdnaqdhehRY4GGkKAorAga1A6kQK+bPElGgLc7GtG0SXb/WPe6El4Of2KGkj0R
kxHvS0SwYtaXAgpund1z93Mq9FVWsnWLyZXYI8PgYkqFcIjpHj7VsLtm7xQ5Y2tD
SLE+4HbIgYTE+Myee2NR1qG4Rq/z6mL3QazFu9Jww9dKYyON0rGzSm+SGcTVCqLt
YT1gBdSqOqEi/AN4I45gBWJe6a15ix3TkY5iSjjHj/NLnYUdN3Z1iFUAe9lgrMfr
Pyqv+EhcNjONyJcsjeI72aPgMJ6qKwU7IZz9eufg7jR20mxlWXIEp4OkiuUEdUvg
+mSbetFseF0CGKVYwzEnAg==

`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 15312)
`pragma protect data_block
DwT76pIpyqDxkiNVXmo5psC9kPE4qtUQ4KTMpeSIkX37dsiLQXIYd+lYdgl2yRps
VKVq/xi0G+9P0+0xaxJeG5a4EHMxYvY+LqjcYmMSXxo/XU6bq1vhFb02olzDegao
E1I1BOzwYsoTJxBcpWUOF0LZ6DFhW/dCAZVIt199zlq1v//vSP0JmQ9QxIxicLl7
US3WaJ8GiwOLb1i95JBbLLjk+yQwROcwy/W3eKMkLyO38m9bqcrxCiNTalT5pvVT
omMNxL98RrZOIpRDFNBuds49Nb+UR3epC+nJ1s1CousrZoqA17AZNmd/wmPP6Syn
Rncmy+DDNsqKTJnMmLd8pozZuG+onGOCenN96gwski+jDtzLSHEfC+SyoZdH7y6S
ZUJTyrSwOwI5Yf6Z/XUcdNV23kr7fuV43cQLexGuWaLVei9OjJwY+WP7JhdX1/g/
PKHsaT957OKKVNmzpJpdqicQnYiapQMslLT07yyKE2lhy6e+zleseH30DgEemcmL
h2c7fzURNos+v5PBVemz4ZJbjVUH7ZmosGKvSUO4Y+GSlcUSX9nMLwo2SNYB+W+2
/uRRRRCiGt2PGA+YDyP5FnJvOtqWwTBk/yf0LdgRvB7w5LY27d/d27s6b24o+LXL
sFQuySR9zhIx80I8rfe8LGWkF+lE0Q7U+cC++byzI5N9MaeoJpDxVIq9coyRyDa6
49nnn2V3/eXrPVx68uUv35UEyFHdgH5w5fHhKwoKRWKlsm4O3DPxuxiZUoIerMF8
SdjlCzBPYyTqJUUy0eBdM1xITzLBCkbN+KqOS+UQkdhl4J+foqAVq6+mByta0Trh
H+jba+491uGZjbTXsmxioe7VMj0IdtrNWP1jhvbFnRChAmj/+m9QBG6rQFpQQMYt
jSRtBCUpFuxDSZ12d9TvakWWzQH+du/kscc+dH4zxkOczg00frdHmvYVK1MwGmwb
hoqXgqPQe68ipUycAnbiyFBvIrROjAsE+BW3E43YfoHCDE1jeIHqD7ZfpUhlvA1f
WMUlxypHqQ3viZAO0Nq7wV2GeZ4GkcXCYiPUxjtNBNDxltXQyQKTOYaxp+4OF9Ri
4OsrnIMP6ZjQOt6IN3OW9GmDXFMi5fQ7pTjaE6BeYW7E4VY93n6VCESoPFbG2bWY
XCZEPsNhyaWzSc7/zRiABdl1uY0htXlOMKJLjIkzaV8SIfQPM2FqPt4ziAwBegKP
3kegp/p9qxSQ1TgN1zWNF+rihMZvvYHOm3y01BaEOnZ3ToGW0O6ZWoKfI7BrnuL2
Pv2VFC+q9R0KL6U/sMDDUMrwEm7A5ugFsF9XfxtaOX6wYrYrWJR5ToN3PXVpgRA+
dnBz27EMubmmxMtpPIJkcHgtjHwdIrnYkZFJdoOeJkfnqzVDA4m3N5VLOgKuEPIX
Vb6ShX4DXVdMGfcXJYUHqvDDp0IZLKfQbO4w7ExG+TceFHvHw5eoFD4aA5bTVAzE
Tn2sEZtN20FrDI2M4TS+zZtjmq1edMC8Q2JteNTgSwsg/X3h6ktOEbQe6ckuAWun
UljyUNQVWWoYglXz2qarUjxiGVPDqLP5hB8G9phlsx5kZaowKf+jAuh18Wt/kF7x
nwjSf4j4LhoYAdRpGVwacJ8crl0B+e6YIZ8+BBFM3hxo0FpuFMgSLWh1vTcc5QWy
4uk3eYZqkelcxJVVJGOoxGHqpbwkb5T8FSwnDGCXka1Z4QetCK14SqHQrdmD1gi3
02ZKdBmhakio3ixT8/fuHQ5vtbW1uzT5I5sF2W+YKA82Qhx9Ewb3Htviu8OXKFnR
FMsFgWi7sJrn4FOOp12Aa8Eggs2yBvxodb/YEKR6R+P2qvNEjU50q0zcK+1Cvf9E
j3SPrGxyAApO0xyuo4Fj5WwfefVCeFZcOSZ1X87JpHAoq9uF+tsFPyAoFxo+j+fG
4TGxLJLAH6cpDZ72qu6m5+RFRL32Kc3XRvpmlMgnf/sXaBQojglG7+WTv+clLfEP
zn7+dAJPgau6JtTzE3h1Bs9pTeZw8UAuhlYBVWUviRKnE7vhHqMSdUKPSXujsGcm
2+LPy9QzcBWqOlem0sa7EyCO/Ly4a7knAbBlihuyYEWONOPcdM6URCNZWeUm7Szp
HUJkiwFrgusuDRBfWxDZo1gtzTbxX8gwDiQDDp+OPuGJQPNK+LYILu0e+FKTYnQZ
iRvkddVdYkj3gfcPZGHLy4XHCfTGc6C8e39lY75djw/AGEmnokinnxdrNA+5y5JU
yXqT9R9K22EPqLI4J/TcFimDZ6CAl5AuaSmYwP2OVMJzhfDh/rRmaGbuVbwXpdbV
Y3V+m+iFa4wd9yzfFH0loIw0HqcwlYLz371VgM224qdmtgakve4gMDLi7y0gWb5M
o7lMshbXpF2tYGvp/pT2lGWfePU+1C7qnYj7Yxar+y5oaeTOVTxsUdTiZJ/2KQtk
XSyETrYIAMRxmPVRUMGx8Qdc3j8m6VRBrAggP9CurN4GjLbaoLEUTua3TN28xZqO
QofHSttgaSz3hBO2YiPFC6g8Ch/OhglinSPhbUyocJW8ob+jF/aIWYMN29uk7Hh4
/ZfVMDMx9rGOjY9+WWDLjiClAu0VS89ENBVV45hYrboFWmE7YFt+7QzUVaXLaRQv
qV+SsPU9m/TfEhcqFTjfTtc326JezOds8v/uHojnMWhXS9X4CfBKkLS12EDXN+h5
yHxYDn4IkcLadOPQiPhaUsuWhZB9GbDT4KBFrRx2qHXfM7RN3VajNp1HpvlIEFz3
TV2o4eH+aEb1xA9flXcfYCwazvq447d+q+R/6iECsx8dHzlnDcYlEY8LIhfqM8Jw
k3Ty5II9gzjbCqLbVR280mc++ID19PtFcb8uc5qnqyACPd+/wgNP3mewS1oEn+Ik
7FrAU+NMRLoACDkxIp55+ewgAWvoK6pD6eqNz9upS7EkZZt7VxSeMUO32VFNg693
WLg9Ud9imhOiA1KAI0zNrJdq4Zm3uoC60VC4LJiAQqRaNA8RlHESZy5PbviQCRd4
vVzrTt+LwHIHdyKkDSnhlz++h7cVFrXYAHugHMoSoyVXdrSrjI1JfJw32Ujz8a2k
BzgYXVQ4jTndz3zFxq8qiizwhcU3JspzRtRFsCVxSapAZrd8mbSqBgmZaKuCZTX1
8j/2I8AM4uWg3Q/l1HULV+kGja4w4EuS0mzHp+7oo/UteQ8xgle49sgWn/QumtKm
AVe5AKdopstmX0gtktN6PIn5J2cckWQ+hBGlTUtj2AL1wexQujF+Kc/fJzPkri42
BrhtE+CKvBF63jgGoq0Vy43E6E6yaTVldw5cSP7bYXi/vQEO2ONDD0MUCeQPiI2B
5q9J999oh+pXrG6XCVxC7Vdhob7ij/vknHhEvN0Uh3EPAAuVGnV5d+Kb2ys0Xa/C
F/94USc3kjNxRbG3QmJ5BmfoFo93QkEDPx+NNyfn5RLu1v5t1fmK0pPgGhizGbFd
h77e5DRCwX5Djtw6+OnmlLLSRyp+XV336wyqmyixEeA2GIFWxMqgRIo/12IMLFJO
5ZtijfNAm0W4lcU0epfr3K2KyUx7mgGW46afK5bLl4KtiawziVCND8H/ucMB2Soi
MqaFSi/K4rj+mJMQVbFv0VRUsUI3EHkYpnXuCVYpPN9SUPcUWYGDM5f0oia0P2Jf
nEEX+Fkm55LSllO5I/Eb+MlMxM0OQPHBPbEdsGstFmIuarCHmNfaDrXr7kflZ7Bh
NFghEJ/m2rWNHAFpUbKWAnxPo3cVG3kcYgfxhs/WfHTV7zA3evY9I/xMO7vl5jE1
K39FvcPVtAwKzC9QZ6nhF0GJYpjJ6vBSwDufqe9TMZKJO5L4RW+T8nEQT6uNn6Mj
NcYHQFrreUorOFjo9bUvZ4Gpn8T+uBsVhJAtCQopQizt57Xsx9myja+LYCmLNstL
W2YB2XADuB2FVky5UaRs5ZiSiO7GY2Q1WMiJngdIKgvwcZVisG37CXjsBdNLE0Dr
Ycgl9DxqDudhEuoXFfaThQnAJM3gbSQ3szePOFd1Krc2jH/XCrQVUQvuQ4XItN7Y
z3eiWI1CconkzVNClIY5ULqQlqGlCEhufFe5oI4qwG/CKomaxGgIK0Lzbn5H449x
n1t0D1pmBivzhYwcCtNkqYSrw0gVvHxDJMSNsScbZL2E9CIcsbwIWwvaqTTp42/k
mWoQEdoePXmUqmaNQbnTYC9a9ksGYSFSOe+5O7sq5SfTiUpIQm8kp//cWD4CcnHI
23ai6LPCluVRtRcGjWi47zrI5oa0WkV/dj1Sibuvw6AQEZX9kb5ynlF2Si56K0/F
D512GUgE1DiHM0+2IKlOJjzZV0PMlB4r8gqvDX7sCuaBAwtzAhS8zrrsSr28KVsl
peDyUAeNobCTMlwW/lrIPC5tZSnyfM4b8yscFgD6xvohx/XS+FA4/uaxOuO/f98L
j4GN25ORe8Xkx002VOjJwiuVc6PBjsDVcd98XXgJ1B9bsH8K+YWADD6LWMN79PD3
o7vwjLG1RQBQ2J3QgeXXC5GvkHxcAlUssEKOP0hGvymlc5squl7tOb95zIiawP3V
Uf6+cfnXvpHeTR4fDusotQoowLuqtOtKixwt2ajlztWeROllgYAMbD8VBLh2CBFb
Fqv+duViAkRgqJyf61kJAdnaIbZ+62XcGKp5D8Dj0PC1CunujlXALMKtuNKX3Ak9
Rc1BbE1pT/K8FWsEd9TXqyxd3iv139SqoxvHeDzX89iRzlPSHqpF23IeqQrpMR3+
pJuZlpxDwgmkLnaKFOodFJYYWgBQ2J1LoFPezvGkfp4kPrWGiEfaEqrRfO7+IMCN
98Tb0IjnCsb79shLsmGukPqC5ClB5GR2JJBtZN1KBZfdmjJ7QzSSESBiPUQ1EMa7
5cKfv8zDVGtVLkJooxdphP4/iyCL6nHpN2ZObVl0xOUATlraZPTiQh/QDAHwwRLO
ne3CkxfjO5MCHifkLHuKBCIn0U6Qln5VO9PBRRGKpkQotgWBi7shcaCMBAeoc9+p
w6HhVNk6Ddc/3tk5Bs/Ts1wW2UDnOGXxRH0HylMtM891T5wtE7cjBtQxYJ8ArhTL
9y5SdOGbi9Pr1Zt6mO7h1heeZesMNcAxbDAEIJi5VYJJfKW8RVp/jkuRY6XtR+Jw
jsRo8vFgO143yhCmRhy9woNA7U8fz3xqlRj5wICTctp7GbCSql+YW43+dgnEin05
q0Rl6ZWhvC88b0R4ueJoQK/NOCdKEC6+kSfHL9GDvAuCny5hT8Phzz7ZaL+IGqPa
4ahIs96mmOlN3CRTZeKZbdHgyyT3P7OW6yDSuKQ0AX9OfuovZoxz4DYNIK0bDvk3
Qn+gh+BFbvTdO+vH1/kZu6GMJTe6RFL7kc54q1/fug94JzwqjGcL3iXeSpFcJO2i
7LNXxdYeJdtrNA+9j46OsHpnUGanlWco9JyJKxG74FJ8kHAaMdSstrql/yBNVOV2
coOpf1llaaAmnNdiXSiLLDo2z0AxoT7BDHKM7DESi4SyYLQ/8Gvj/KhTPvySpsA2
I4EHZUa6w0FqniltGuE4yRfSgdPKRGAxn9ZuMH5HYqeEIe3vYJZ6hcWioNJ3l/nZ
2ekfJns4Vgtie96qMp/WDcDSnnHu907WodgBdVWKxttwl4Kg65URc1+PqJH9sdJM
67jef2BctvsEG3T3j27+79R9XKOiDfYn0RFjqHOc1AUh63qR8JZ8fkpEVtGQuK/n
lPUKIeTcs231Do5T6KoVP9Ghu8hmbMiWOFYzkgjgbrb7tOIheVp6PV4MEdvz10T2
or6EKHZhm/EKOuYaTOYpnUDSQgFx9318afw0e6Wkr67A58zfJzYHAW1//rzb/0gC
V3ppeFYhdZz8Hcec4SEX7bTdAmfulIhaXguGl89eknMCg9Ic2X2Eripc1epP6xdp
JUz5nd2ONU2ThjMqAxjBt2EmUA+xlbs7i54pJi7Am0rHdLP0dzshOAESS8jSyLrF
gpNIv7JvLvRFFEr6snH6j288ry8fCt6yLN8mIWjk0pHbxSr2oRHBFQH2ppZu1Gj4
LxBaTfmM4s7EAGC31qLybWhhyGclP2Pn6OD+yQgsy2shpBUgArBbF+7nROCZlgAY
pWhvA0CUN1lFLNtW6V9UUO0R5cGztbneaGYc04rpTFVM/rrxR0h3x/Tu1PWMopGR
qQ9MJgq8r+l4S6mSs/zkGp7F4oZD6Fbvnrc57r6udUppovWfGYATIr6vsHYbFiP5
K3Nk4vSw5L5UonPtIg8LT1y7zj9GCu/NWE7Yoiuemvq9F07Out2TPEP5MxcKZLFi
TkisK/EEmQlcKJtzv0o8L3PKVFRBfO61oSIcvI/5Uweb9rfUL5BQ86gttoHLBIwn
u2xS7kOFpsGRfBYkmFWJ9JzMpFb8b31xzmAmZBWC8ph2iax5lRJ0sTssn8YYDhgp
hgZhgTrawWbtTUT7jIWUxKBshBx3iZ1WaCBU0AiJeUoEiOx5XjDrEBeokldC286V
VN8EFOVhS+eyONrNt2nOcVgdCPfeE7zL5AsxhaNF+KgRM77VwWIZaCEFcTweSTi5
Hz1x3S4lFU2vSsBUMEMBn5/idRXWrvRP1F4RaLupgLu27Uiw+jFFIrh6DbdVfEJs
auY829FjaZzOt4Z34p7/hlRFkWsqvy0yhXpyplClXGJRO9QC/7bT+wOIhYcwaPkY
3XQlgRSKNivfop93X9Q+RfdHsIwepkZHKYZy2UsfOuo90BDnLHCjzNm6fR+WjxIx
gtYoxo3uY4x35MsfiDbnRXoVwpY3K3fC6oDdh3bUX6k2eiH0Qdb1s+rzazIadzze
hCCWuWwvNXgCpAkb29sodZrnWuB1FDgyrnLqyMDvvta8dirh83fyXt9RAi7vwyX3
XkRSphqsIGFRA/S6dYcEBdaZnZXBqqEHyvhy7b0gGa7nzZQnbjCDnpYARtqv1QSz
83/ewYUh3WoVyTdk1Ffg/xpIglObi66Nei3MqxifYIaGPYq2VKOckKalWeYCtTCB
8M++MTFcCDRFYdJS5fgUhkAJuoMM+nyVUazWAei5yuU89DQZQlKazizcHszYb1xW
1DpkMAO1QayJhpG8Z5RXphV80k0XoMfP8GVyjeKYkfSiJ5uC9DOOxoBGCpCWsIf/
hfvG//eNOgHWhWdOG69rvhwDOzvJ+MmOdf60+c4ujA+FrCPIxTdNEBbopvJzAAC7
6TsPqFXZ7Q5cm4Rcyz4mKmsI3wS63oGF2+O2dfMtD4dbODjU5YAPJnDFziPzDtfY
cDFMfx3BCzlzm9iQpwN44WVa51pTjV8g0YnRKC2P6VHYZDjzynZ2C5EX+gxhCkSY
mPJNaOPbW/JnLQ8Ttjpru4pUuBhZv62nL6OzNI7xss/j9nQYLwOq48piwk7erujo
H6qIefdmlF+okVsyrY8yaH/dN5lDhKVVY0ufIcHVfWL+2f1ravRVShf3mluJ9FLT
3WZJ31hrDEhwpJWjBB7W2jz2M0oXrMh2mqMAPQwticR32mDpSxh6urMGO0mPcFaM
Lz/DZYvgDKPqJYiMCzuAjDn2mV4nZdRi/ncnHPuqQZ9OjCdeOIiFf30wDIJKZubJ
D0ts81d/lsbaoflOkNYcBFQyU6zDgip+WrX7+R+4N/0Q1sa2/HOcNrwfh2XCd5K7
S2nsmt2h2e36bOfA/6Yf5RgSdu7hf4O2KkojJu1SQGIcjgzTuLDIVukoejrBX+lo
JPzzIndXMiLn9KFHqKEPm3blgFbD62a1PqEbOTPyES/oseTQv3SVi7vmcgSm0RMF
YgzSXUudja/xb9KyFJ8vUrUe8PM+u/Wpy5uhAGoVRzaSyo2pyo2VKiQ+giyyG3Pd
sfR3Uka6/+zhUJZrP49R7Tb0DK1OdT6M3Xdqd8TJLMeauJGFm+GdLvELoDiNfJRN
8fi28ZpqJoEB7JxA0ej11iC5v56sv9Bdksjdr6HACFy4VpJb9d2hYdaFSs3t7njm
26oHORQyT3plpbWQsWvuF9Q3aWBVxNnY8CArXMJUDMhkrWQngMR/P9NPlw4/ZYOb
e3klJyBVb2b7JKVvetDb5CCbZVabaTz+3xSNLJST8LJ5MJUvHf2yrHdZXQTk5xPw
jvMo6CBcCtUXjHvk2XHXWkC6ec61VSKYPK4q+G8D3z3DlubT2HKW9oflglc8WEEw
i2Eum0YxZB/fDYREn21BDGAa7Sxlp0NYNFqLWDTty+U937cf6zWiU76Bh2M9kjv8
1ulFpXJC01LaNBj185vUimWZtqABj3M6vUuoTx6sqcmj1EN0s42CTMITBAwS6Qbl
KKrDv3rm9HGMTvf2LC3AGkpOE4SPARE70kviHLSldJxAjo09cL3Lj36wozjvBREw
LbFXAWkt8kmuF6a4DKBIabWWle1R3BI9RWvVgKgab0teCk3hsLTr0aYl4mB0uHS8
YeHZPLqJs/N7/28rihlR2/1fs8z8aemYrf3ZXnyTsqhVJxFWSVv3oVExcjwWmXEK
OTQp15xURtVuKFPRyb7YY3pxFtw6bAl/PgsKIP7NBIdrvHdbbmN9tW4G2+k00L1s
GtLQA9/DPZ241kHpYEAO2qj9ayqb0hG4TROCzOyI9lRkmcOnNW14AQiS9ZW2VuLe
KbKd8TeYWtao2aTHAN5cQwFj6RaU6u5yUT6uRvhvR0poATs76MQNJsJNibNcwK5R
jENM0Uvbk1dVdxadyK4O1lojgb18NEtYbT7Aywh08M5uidBJhf0JOxTGi/pH6RBX
ouBzh33j6ox9i/y5HS0ArBrQBRGElLKIwX/uddsjBF/+djxzT6u0KN2iAkZXcbia
eNN390r9oKsLEJA9PAi+0f198/wuhzb+qs/EH+p2loU2LCa3JLNlnrlFr4GU8sIk
ST2a5x3CDZNz1LV5H8kjhw/ZbCfifm5GgM6aqg3KeaYTsWFyUTIAIe8w5bSKMAk0
SQFCI/Wb2K0qGTLrW56ivewzPz/HWcTuD2SrEXlh07JW23nhiVbvaUTP4lEcRmvB
EI36d/jgSgCbRn+KqGm6fn2157ZdQJ61pE8k7/hny2ZRa3Ul3p2aApuStMAgG9lt
OPzsPj1VW+ywND0P6SAkPR+UL3y9q290BSY4FtyhTpZ+T+MPV3PdzkLNG47DuQPi
Zv1TsgL61lbK0O+BBblDRRO2IVPZSe/MbYAODv1Spu1eUbXtm2tjrb62ZiuIr4th
dF8hbIkQF5WN/QTkw6gqRFy+vXK0riBkt1l7cWD0U6BykykPAacNteph8rLtjwP9
7BG6X4vfsEQ1gNhiKOB70iu84k+AUbYvfmpc/uDxrGWOhxEucWv/RKwp7k7PCtbM
R9hSBHNtQrbeyuNem31gU33M3hn5HBuPlaMhbzgPWJa0JNZdf07wEI7xm65LoeOJ
CdkPpruS/duWKKLNzB8xh6C2Y6Z6O2SU2BFU50pOVl+Z5oQ/XGxxC2ItOCz6gVd9
YsaqTW9e9MDy9F1XTKFwD9qxCV7piiR/e0CBVzYRpZ3/wRxL9H/IfVp20iSto22d
IhaCyq5ydEzmUiWeRSJNYtKYssYK/f2WxtZUGQN81WXRmzRLxI9TeVEugOucUaYo
GtZmrbzBxRFgjmwNUNnP9f/x54kWrhWsbPZRPMlA96laiFAeIxqOAg5Xv5T39GiA
LgYmDDPfwoOn8jiNv/OtQWh4cejMHe6AzAADXVlIezWijM/XL5iDgoOEcxxQkapJ
QSCuQMQyHh6m3ph7rp9Acfx/HY8MTm94A07gtidryWiursBH84XNySxLn0hmxcTC
N1nFufV9ltS2Ujqzc4mHqG5F4AMJQ5jRaoqVrteVxhP0crp/gBqh1GeDEqFHVoej
K06ezULSES/ZH+SOhUn2avyEMGghGTGCxVa2BUlGR15/+OjxX+/WbEeXOJzIyDFw
qTaHdBdzgWhmOdwjQoi27DIcq0x2Q4ShqbIcPQ/Y+FZSd70Vfn3Er1Uy2qgGoRKz
wkQGDdKJn+kkSjsAYiRt9l65Kml7eTGq+x4gyPej9g0ZLkUTCpjCLarqC4Drzhsy
AjqT5SNbtkP+6CnnFLYTH2Oln2aSEjxiqA7+tw5miRtvS5SajgqtIBWKbAVuySK5
NbFdtDtHxUtLi9YH2oG4YQypNxi+iGyc1g3UELbGpK21wUxsaT60BJcS008+lywd
CIgxwRHG3G9TD0LK14KMAppkGg6yH0cBNT+p2NIvAvmVoPD5JQvmtD1q/RIfXgcc
Lys1Vz3FZmXsgGOPzuwOltKbizFusF3A7C64HupT71njb1ZaSpkjB7+OV43OtFQg
/iTRnAfFj9AG8HfWILXYSlVoqTfhv0GgMn/llgPiPeYPjRXMSl060EiAAnqbowZe
FqFvZu2ZwPyGYlac4IW55hAnL04nffKb11pqSw9a5vpwibG/8BKAP8McI2xlxQyF
+BGQoabdFgmHAra/uiocPQQNwMy8d/Fnz5hq47xwy/psiEYVUp4NAeYW152dxoje
gZG2ruwXrnNCzhEuhSGLmXGd+Xy6RnCsNg0vU00/XemI3TojFS7ehLFe4PGn31ML
Mqr594L5DQSQpNr3iyKSaRbL4tnhevemgyNvhDMSqdAh7eE+yC28HrJ8ouqHP178
skogXXBegjE1q+zZ6R50horIeusXMMh/4Q3KZj+EEG7BnGGHvWbDPgepAMae8woB
MRiRnPJANe5HXMwnu1C6PlFTLhmeWYNi/PUz1ooQbPjsdcxGCi3KsnPWg1IbvZq3
t6WjJhuS7+dkMdz2KSURZ3nZCkToC/U0qHeyw0xnM/PYTGIiLTnqB45ggWkmDuLN
Tu6KagcFU89oK6t15ZPD1RXdvIsVGcl0UCnT7cTLVTRAfYY5m9qRCBnDeOjw28ju
DKGrdYNBx6XlJIyfZijJPm/8av1GcOICxMn1HhqCPtT0Kwh2vF6psJ7BW5UJG4n3
kipuM9twEEBXlIHKv0inLzZnTk/8nz55to2ek/MEZA1zC8xRkTkcNc9s+Emt1MGt
q0JyXB/rV6LxSlbAhp17hI2ZvRxuHTUUXc1FgsxAIfY2KTgMCxEisoR4QUop9cHc
Muq2ncfpNvvwnPB1najeRZ/0UC7nPV016fZ7wd3jFoczV9gJedgrNIvJDq6ZP5MG
0h96tUBQuWa0qCXv11mxjrwZeyB2rVIM0SpueZ2TtptIMrTgcPpRJdctMpiwBjNe
Lti3fvhtlweoj0XpORJcVHlAy47cFvmn6tQvONjEhiNBEt6iRm/V7+yZ/yLdDNLz
NgsbqyFs/sM0D+N6b6y7f2TC8uJSDaGz5ezq7BxCRcLfdDef/4pCAkl/Rraxj6HF
hXX+zj63Yy6hPhhivtnd4qGQoqJpHXPAF+KkcxgEfbgJsmsVMJy0q0vISZgDrCgw
5wMBzoWJRlLLa8/GD1AZjjCfU3P3THvYoE3N69EfuyniDlzSj/V7TrYBDiILQ6BT
TO54jQ302cfcq+tKzZCpOkeEoyhGWFuc6zfDjhrUwJ5eSnse6FCZh5QSGPc9tBih
AFCPAC46OekNETX1eV8wPR7Fn6pxcGyac56uZkKOY234X7hDNjJfggLoRsfr+Q4D
7scWPZQVjPlwgrQk5AKDKMPbKokPaLRKwzT0d/SOm4Nbzdbk8ZF+u74KI2W2hU6d
+10jQBnIxLuxRxl1/6Y1gC/7MFiOX4o0K5NZaVLXqE7IzJlqRPTnmcnR5tNcXPOs
M+he+k7uAQ+zHsS9Rg08SQsr0LwV3KS2tyPHGO/GPDwYxEPmyYAZXbUcHkXRyXxH
h0xPWltw/3lkldeA7PxUj8AO5R9c0OIRkixsf3O0do8wJIlAroQQ3YpyeqiUEZze
3gwI+a7Mbyv6cI5RXfngGJRBTIc6jMkItmSr4l8WY+2qJ4QnUwu9cuThT0o/ySBQ
XZp9cHK81rORxwAWbfG7tmqqhdphMyFrZLSimD4doa5iRVVLDpMyl+aF8dK+UiBf
AK7p+3ywyejmSmivEJ3AW4bW5NTxwiDyvpZODfKMlSFSs/JiSIBiMcXeTleIWtag
zUPKxWbP9BzKasvFNGmG1fWtpNHza3VMmDeJz0ra+76/h4VzTrUmJ2hw8/+OYTwv
HrJtVTN4YQiqdo47S9lGd+PzlnAmXp8+G1pIev8tVu8IKm/Y6fBluuaOwrYmJG/z
6y/gPgd00/REQtTiOl82Ka4P0kLwVmWyyQ7xQONjI0mhvSr8yFu3+ex2cLsJt89v
+ebwBg/c5krbb3rW2FzJh6uWO3dRxaDjno8Ht8uagjjUPqnxv3RMCVYA2B95edhT
zIZ5kIQGtNLNfbQoIDBgeT2nc7xI7LsTisYalCPF1ChhYeOfdvjsNibWzoFQ7F1b
HJhqNjl/Z/x23sUMZW0YYkzQFla5zQFXTRZSqJsPuB9h9mHqHJC6O+0BnKZj6Kdc
Wn2iC3cuVIncWNLAiJQUlYK19guqdwaJq6T/Qbqs8LrzO5cOeJNUU/NKy1+AZUIu
KQ+/FvWtmE3xcH0IV8YRAUpcvXfARBbEViWHr24aA4N+x/ML2YX8DWFJqUlfJXqa
Jrgoci97mYoJC6szeWgsBLpYoV2o/Gib8OFzZ/JcqF+5zTLcatv9Bz6SeKSnKs8o
Fc+b+OmSx2VaO94Lq5O6p5yCWS+L2yVvRv/7sv6uMvt2wYNrgHmYWKAgl2zriU2W
2EmhVfd0xsHrAlTeen7mI8s/v4Sdt11GuTaLdaDds7MOR5HjLV94iOrY7T/wbfv1
IV4qk1hjPCXJJ5RrH37YE5s9Uqt7Jd125HRsoKpGYrIiREw0fx9lIIgbtMLjjcCw
uHPQ+3IicVvtKg3wIOLkdAhvEhe2Gfopy8fQV2MPcDD/cpCzqSTjnWW12f93sWcC
LnaFsikv2vZXuKUr73BI9BI3Es9VYDW7aOwt3e9gzbSTSlEiehYsZsaY4OTXlE38
oSpMEozclL8AQduX4IIibjyZOPFfVZ+43bun4MbMidf/dq11ZNwiz7JUvHTIYcxh
ymOJuCluX8yCsvMf6fACybdnP7bDQ+NBxJfuoic4It0fmKPW1hmgIcD269WAN7Hm
JOptdoNIwY7tBkviu7HHKEqmhyvzc92ZsxNCHXn1nTzlgG+3B450yrbZwACpo1Wz
3TfMnefvivAwoL9nqlg1czpoJFksY24bxd6WkzQl5LEXcqJpHPlCRrhZqqbK3V9+
NOOTDQcl4dG77pi0PWOP8eiNIFH5mGVXMCKUIYHhezHz4LYMLVLXDnp/sx2+wnVL
hZURTpQYgo8KdBrsjUER8wTeFqPa1xZj3k/soRQgxljQfOHgMmXlY/L8k7HS6bDQ
ZFQzqxGfWtUjXySIpBBY02DpfvLWkcPnXJNKyNH9QPMrNxxV6FosIYw+7BTQYnug
XfbT5sRgUoa6oYbngIX6+N7t/OYXPsleukK8hQls9UsrJf6wTZu7WMYWEq/6hAsJ
mvCo5r/wnXbMa+Ge74as8Nst91p9mYOl0/IXP682+leIEuOtvRd+nQy5P4CVlkji
9zy2N40Jj12JxBDEC86pdddSXu+w971nw8XsmdgFYe1RkxqSt/bwMYjYFvVxlciC
hkB31xUyyDfsp0FJVvY4NEHASvpHqAJwf5AtT8As7Qcl0sHnyljrsOHkk7/Xsh7y
7YOlaI4BI1RkS81kY1pHbnbVb0e8k3VBEsAqxyzUursUuHAJIfFDhyG2Hf/dYtz0
Rggvvvvgryt+VReBxDI1vFAsJtHoHrAhEijI150RU/5HidP/q51KeooIaGSQxwSI
eJJpJBO+BVwIerz9qer1yMyMcbQSj72CraTRtkmFHNX9BrvOGOV0m7izNqwff5Fx
uviyYvZxnT1YR68kJr7QyIAxeRIAteouNbsJpXN3ED2Azur2BBGueSE7A0ntf32n
2cIesYZdgz1eiO199ceO67cwGFunA0t8XVmV3MLH3vC2duIUoaeB0qkZlclPn7kq
XhiGO9ZitCHtOxqb6BlWJAsZq26xMmJmtiQBONhSZnX2JlaRna5Ux9RkKz+T04v4
GEXL5ENwR3WMKrv2Gnw+oEqYIF4rmaK5BpUHHEPxmrYPhxHndaG9/zuWILnst+H3
sBjGAURebmKdpTk+PECEFKLWv+gxUThBhjRmuBBkDBYuU3jP4ltkVU3ZjFZNwqaV
4GMhhu9fLICJJX11JFH7CwwvTt6NBMzQaNJNzoj/zaSjeFljKXWZtZc5j6t0h99u
OkTaPXIZsmleuzMs5V+S6zbLhZnaMIvFkQN+dlXxh3Gt+WDrv5Ja/WgXAYSp2UFp
s7f5Y0if3XRx+kGBUUCJZguiS62H6tA98j1wzOuioKHcxLeXELfWbTGeDc4l0qjJ
HJbtchpFluX4yKW31aeWQPvT8TYhPBkLVPL12J7upeXxleQHduSxkyIMd/lhiXvi
VbGqEoksw2SbLSxlLIqz1995ZK8VO0gRFEj3CL9HCFLdj7qpDSCX0ZGwHAzjP1Fd
gW8aEiKlfpzI4+xd3z7BBM3vLzl6OnWuKvL/PA42Ta4FOpMnd1zf0h6EWlQZQs+Q
GLeOoSADQHgZnVZP9/1u+HUYM5SA2QDzr2x2NRQg89Dk19cR82mHiVXgfVhTG/Nq
K6QKTZL25ejWOh/D8Nm1rvEuGJhtt2ThRtOo8NtW8KmMxNNqtTHIy47cdtNo08D2
QJnCRkL4MQE8v9DpVx1WnvNLgs18EymdiDacAyqnrjWZZZjkAIcrEaKomCi8jtfw
uqOJMLoNWDg0bTNe0hib87DSUy2MypMXcjoBsMuoSFZPae6COzD/3rfWXLWXM8Qg
Fa2Up8xVCl4sHFn9z4BLOqYmdqaeBij1+NBsz+4R9yJeL/aX02Bhds+py4Y0XuFb
z4GqX8Jti2r1CPsuffobbRQFt3G1WqZZ0IcCEkwgEY6JucXGRdFcdfXf7qz5B14g
1elJ3UoXLn5xvobq+3AXAZsKyxffjGce6SUflTTqxftp8ZZmXn+mEwAI8C9ip2bJ
N0024TDSjsAd3i6pqoJtvmNaeXUmNvFJE3QH5G1J1+N+OngOF7QHoZsg1q2vqRBA
jLT0uEZu2PZCxdzt787Hu5pEobqxApHs7jHqyGkK/gxK/OmlkkRIdFzHCzbVH3q7
9YZJIbU9YAf/mmLZtD8KcBhLIzyV3ul28eHWVaw/LCWWFX/1UW70yBonhT37jmQo
QUg4ndDWe7bvJyd9ZOpG6Pz9w0wt60Uy734Vyujl/IufL/5t+bnIxcEjkqW3fasY
LD9cefH6K67AbTyx5GZiLkteFhYLPN8zWsB+KTRwTKZPFeSTrgeZaCWQ0muWU5ig
euPNf9bohIARnUzMHk2gu0BpqraWN0/UIKrADN8z7Jy6U/Fhq60P2iBr+VRbl4JQ
Wln/NaQCr29DAY24op5mC3z0fPh64EjDrxiGa2lwPTf8JTWNb3DBdLGye0qtxrLu
L3okUrUmYZjGfMozafWigUSipoRbhMuM8eRTt7iOmLhzBrPSYyXWDPCON2pzftDa
pBBwFEirI16JHQc8G8F1FYIIyK8ZxyboyBOlAbZnnRQ77Aft1cIghe2eGXglHKjV
D42iUox6UsUhLnxTcoc3iq0NBjOAwsBS+EmtENZf+f4hP3KT+9BuwSnX609ckCpk
gw3Chybkyqu0Wos1HINc5+idmZmEqcWoW7k6kmRAylCMkhkF/tZTDzYh9yd0VWAN
g2GbkDQvJw0TNYasLRm+VdIJ83ZmG8KVC8EuKaWhaFQbgxxxStEayM00ugH6ntAt
bkD6Q6ael2FkAqhxj3Nce9Zriq4xFJXPbU67hLf2xB3rnvPznD2tcKg/XHNytmaL
g1YfMuTvTco1lDD/wZQ2SMsZXdTf8Ow8b9bM/q88sZTd3ahHetuglcbrvZu8+MfU
3OBZUQH+JRf5wDPSdi3Dg2qHm/qmiNbJtuLS+I+WjrPFnge1MFF/bR+5yWHfhf6/
XwKfToYmzsiMuc/g1UDqqzO9OfjWS1MwKuuqLbBERB4qVEw9GvYrUWNC4UroJBU5
qtL/hZrw4DG1qNpbO8/VStkTSycXTNK/9UcwKZP1rVA5wQB83IQR7fn7Ln6mgnfp
77tFACK2/lq6urqJcc4ULpzLIyCmFuiB8hGmPNg7tsnhiJ4l464zT2ZPfzSvUwIb
a2HcaFJI3xQAEsvN90uEa18J00ayMJUrpSVgXDVEPqfcuQqOEXK3xuOjpUlm/nI7
qhTiX8IzNtubZ+NEtFCQIBCqkht01H7hRsD7j73lWLdSclif7wUqcgDltcGrKNj8
9lF3zVoRWXe0jb2jYKUZysUYoGUDCYCx+E+s2i1SwxEvLO0xDZ/zJtD2dg3lo+wz
r9pAcvJyhRJvvxX+xco2OfzUHr69Tv0894+r1dI3s78Gq5mUMR6rVcAzqzT8Bdze
WM13PEzZo1OuL8+/5coycxZEAlDlo6CHQKxup9/O3La4+LxMe52ktNa0iy8WKtwS
KQ52FaJTBVwraeDaJ8Vz6OVNP85gFlXdCnNMSPDMTgtskFNWYSIqdBeb/NqaknUM
3MKTBT5oX7vxmhuvyRtZM4BRpwQ/07TaYml0kNVaDHZXJqnZK+aK1SdsjQRo7YJ6
N9gLT4CiP2da8GoAtpcVwt6yHukclZkzEA4oen2cfsZWt+qphLzbpbOvsV8FwECK
y0H0Nz/l5s2W3TLitSI0y28IEJO3sH50KC4muJLKS0Pn/B/9qdTVTiD/0ztNsqBR
hcaEwlo6rIzSvn6aW+fFvGqgxugHqSRRLa6rNoD2Cpktm7ANlKZZmLHkRdFM3yvM
sjwyr33Ut2wh6COj/UUtVIONZkLpRYNX7xVk53V3XKfwb3/PjkIVryKBesndTCbC
/KdYlnIv8G40o89MdV+OmImVz9bSWcITMe6Dkjyx8cJDZxAXtVxIjcm9L/+tfDoN
EXjKLdTd+R9vkhdm9CgKfVQGgiqDmJ4FU/AatbQDylCWzPHsLle8RUxJzNZoDD2V
bgAGQx2VNVGJ4SICCmZcAox0p9EZ4l1hc+bzrjJF7NrOj9V3BOmb7Xx5cmIGDJ0K
TxstqMiij82ReQiEaDgtj34AQo+YwxqcsFoUaYl/H4c2Cl0c1q/f7jAm+LnSYg38
SQxTa7BLb1JS89jCa0J32ovroEeSS2xZfMFjsJGr0LKQvhXShmFjqEpOCoeaWEED
ha3dqc9IunxTeqmtzFvhRmM+P9DaGJ41pS0A94DmJ65aJHbbfml4KWdSmziebf8n
ftB6w2gikJmld6SBGDGOJS0+n3WBrtQa7BtoMrPi2m4tiued9eGXpHanpkSTryCk
OWg5CM9yY+Hp+WJAsfecqIspHxrB6mDcuPdUTFLYlqWm03eDBR8xdOgLKxBapzXs
yZOZ0zFf6GF1horlZz3BQXZZ2ZQk3IT/fCvtGzIjQkF48FQDYtlngUxR9LeSsInz
XEKbHKQVDOtkfbB6w1E4+7KlVUra2WzrhNRmSgcK44qrz/UK5zaAu4rhG5Qozgw6
RqexgwQF5YpWmvnZI7KNh9P2xPyHN6xd+q7gfOtfJWZH9aHFgsErb7F3ZbQ88i47
zxJEmI+xAv46nOxSzUeB/RQHfFFm/fvhSHB8iiqJhisbjeFcCFPgppG8/HuFqOBX
aAXJMOenXIsiIAW8sCOqvG9qpsYYNTHwvFsnxC1Y5YgoSqbV8POdRgYtoauRMhkU
EJK9JkadsdvvZZ46xsmGP3QOP57gvou54Rr3fdHSiCD49rj2ZCIiMZta9EEOfQWU
pmidC/kW3OO1+JjNTxtcwwuitTB08rvtsKmLjyACRbsl/KqpOuyrv7tZ/DE6Ii0K
ci43OQ9/8jkK95ZtYT60OFfjjidMxHipzUW/6NqKyhivMOXGDHJSxHXsM5aPALwr
JnI6fGBumBygww8bj0q3sdQ5dnGisfmpG+NCHtNs9dpUgfbAlib7y3K1nDVNiJTT
v8PRDB55L4HhdZJ7u0cUNlhiVtmwItPOieK5kUl7sU3dAagqVXx9LD0+AMCqEvCL
j9TBL1aKPjZ1bqHTFLBEZQ7GoU6bavXlZ4ewtVIhOs538BStpIsQ+7mnOpIBFerG
IciTLMXrvZzH6h1jn1AxsRSvZ2OB1uE0XBMoVecJhcQbzkTH/0z18ldweIFbOV/K
V3XtMwBuWSAeApvI8jkb3bQoEnCv9y0jM6M5xXrTUFSxSuR5qgPqGeMBhKKBufL7
Mo45Vf/oXwAQ3BPKhEL/xBv1/y85tbKT5BMeWYUhSnBSiND9wy2HSWgTey6u/TB9
EM4S/s2ZPRPrbkOHCoR5XFd35dHQtUwE32WlOEL2P+BsS08VO9TfOD6Jz/PFzmvL
ZFahSO+53O3Ppm6O471duMLzRnwaXL05XoqZYNek9R5xBlQdV+lIpHW0HASrYqco
A6qT0VjQ7e/CpxyUyrl85MxiqXXM6zMrT7c8BWaH24rmQSlS2zROHREuJ3r5dmEc
xYHkkY3HCpkcLe3pzkgIwfGVg5Zf7Q5oAPOaOpWFEityAJomp3gCt3PFpfQOo+qp
NWbWhBvBbiF5H8C3ke3GLqM0EJ6s0W0SyEVTowHqlI6cm+LWJqOLrtQXt3cay9KU
LAWhmuyEj9/+qMkXOpkSmiwbvhwYSogxL08bV78bfYi3OT8WJ2nDm+vqZK+BBYvt
yBXqxX6ANsXH+x8f1pJ4ZGS28OdBTm+j7nKWqw7p4bXXPdDefcUatNEzJ32KU6QW
4ON0U9E+zMaXRSod9AyJYsMOX6Q0fnDp3o4+bDrU5pYVXFnlkH7vmyIm9BIqWHUX
+ZSmTdhYdPZKKar64rvH2ccVR4fFdpq1bF5nFUKQh5IDNW+Qz7yCNQm/ui+dXhtb
bbl8GAdArZbz5jB706rBd5xZMV09Z/s1Zpl/uGp9z9Qd5HvLxyR8LX52SPBbbPro
MG/p+UhFAb8Uz/7hDiC5k4hf/Fys8ym5cZ59avmhcRpZaqUJO1bq84zboEOL2K75
tTUrECfGuoKv4VZr7WCDK5ZCKl8ME8nR3VDzPSX6U6O+5HfxpdvJM3CUISjqWwVT
ucocGYjittZjXemE6fBKFrM3sNCLwHlFNAfdQFjSs78n7yas4BJlr4lpG64zmdT6
FK0TM9MOHOL/hQWMefOfxgqcnXZF/+stAmyC4u9VGH3DvQEtmeHkh2d+k4QnAmlZ
zRZd0jdRr9QuGTFEk+cw0pHGRwz1CqjchSUIdwpo69rphvn+7K+PlddCrUB0oPlO
JLAWpknI118qmMYA2clxbXPKbBAZnPb2SJJylwIF7IdRxZ5m+9aJajeDSsSjGxPD
h99FOXBKyzx0nmdHhYvMiGZtVZgL7C4FlFjWlJnR1qg9UyMUkoGBI9ds7mwTCpEb
bXa5hQ/OgOroxbejwYzzUBUA8sFwD0GYw6286zSJIxcXAcX+TFjIaDM9XkWYK7oc
5ZyaMgBRduQ4Gc2HIBHe2yHlKG5b2ERsUOIeHOnW/UiQGrV6lCpUGnnAEBsACBzp
tK2LA6Gg/LSrtvQ84eMn7XLYE8uOK7uRPZOdV7WlwsG0vpJ5Q6upnr9CuXBct4kD
NRHZiuPXIphcxkwglJV9/cN0c0wgowl3opMOSPyA2OS7m0G2B9NCljAo5Hg620t5
/cUiYA49V3mEMGnFvGB2c4LcQXSk5hY5VbbH3a3V/abphUFbb4GbrrE7v86/RMiD
Mya8ig13fRTk9DgZO5m7YmLD9k5i2KtqHX8+rBkiS9ewqCvqqU7SPJ3dbiZZ3O73
kELsDkSDdgyMWm7RGV/iMHWIO3VuBnwX42dYwTXUUXo4Hu46mXdkkp111JuxQOe4
IIrw4iBwOmms4e+ewm2jZLbFA/9nkI39iBsx7K/ZQiZWQM/k38IFg1iy2TQdtOGp
hxER2ZlgslTpvA/CtFgn/Xg82ywIQ9Y3VlsKOkx8up9yfEXPD1YFm9g1Hdkef5oe
ZD21Nw8kwGHXFbqVNizpthVckf7pFEAAev+Hr9bp+j+ouJYERVZUX6A+jlWY13u2
psYzNDtKP4dhcpKmQRyx8k6mESmtL6PDdevA8fKsKEtVuLW8WVmkObDOlWNWBcg2
NW7SdvXQlzbwH/FXyVDeA4SDGiq76Q9NPmBv0xhnw5MfLB27DmKKjpR4fpeH7UvD
laAGOcqeaTMf+KMmBt9PVzIoSz/CJKEA030rDlcnLHq7nJzEq7ADu+Uie40OwOC1
iDk/rN/VfOKJzXHodN3CHRpg4rSime7yRQzdGTbJdwmeZVQnVyy5WLRzhBwGS7oZ
fkNMEX5i+pxf9b6GeaafKxRPIEUNNH8h3fiYoLYqNJFQZGGXM99ClHzKBh5i9gMM
na0/pEGIm2Tg678aiY8o6eLgIoABEAyCgpacoUmwDzoKFnV1vnhFIwGCSTnOfiM+
cGmasnj3Xhen/b485Q8YA5/uU3AKbyeUoiQgejgkZ58VCEwAucgakYisUleHtoL+
343mwE0Jvp3wLK12kkMXQyAHsosUZBQOYiDixH34foL+0C31wuNxLuUTo2kj6Eok
`pragma protect end_protected
