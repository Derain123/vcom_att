`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="galaxsim"
`pragma protect encrypt_agent_info="https://www.x-epic.com"
`pragma protect key_keyowner="x-epic"
`pragma protect key_keyname="rsa-key1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
VsUG9K4zdGWnTKea6upVJhUJOB2WKHUCJ5k7081uvTgqXhS9KjvqvR9SlSTDlgrl
62+VHwAUqI+UI7NMFngIbf9+KAXw/DEThq4ED0JqIEtp4CR6lPL9RJm51a+aJZQX
bqQoxYoXpkxnRhH/rBNIZIyHwYc2NP7wlcdmQk7M8NtA72QgYP5EnI6mi8ljZcZa
NyTZ1AgbcvtQ/6ObLKtAMlhEQzRinNoU4z+/9Zx8Qa/npkfr4dfecDWUji0Eb+l0
8TvZDjxn72pwT3uAszsZCDQ+718BFOc832l7rF63eEd2YsJFNSCZkQ54gUYvjm9+
PipvfMvyPo6imqnlmG7rEA==
`pragma protect key_keyowner="Xilinx"
`pragma protect key_keyname="xilinxt_2019_02"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
iwPnhX3MMrAzYVFq3/Th3fi+BXOAoKJG0sTCgQaVBQUcnraxfPHFBj6Gba8cUq0L
iUTXrSelXbePi1z5BrEVz7PQTNY9CbdkDaiHnhYiNSpk0c2wtjc4i567xsZTunk9
3CRi9wwGWo1eRepdXHDJShQAv8ohQuQFxovTgT+nFwKtuim5sTMk2G0LuSlCFbfr
WE2k83dHUF9OctVXxWi+xOYKEqBH47NVM/3CoIhxyW9zGWfJcg876wGs7ND6TdNp
dtt3u06HA8Ikn1VaH9HOprODjIUngkDuyEUI3CaA76y72I6VhBfACXs3XfWRMZca
aACdgObFEqZb+AbvfnOY5w==
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`pragma protect key_block
Qfd9L/fUNWcLsBS8SFjylzYqEc5kSz9vYdMzuYUVJP3sW14PYRjQwKo92u4Vui+s
Y1CfTBCJH8jdFngze9+iLhMDkGNk0xxNLlVyP+Z7amVyvrmBmazOh0wBXEllCvZI
t+SagI+xIqozxumQNfoPVm7BRO7MNZ96X0HhFzk7cTs=
`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
qO+0lhTcWx5N7yZ5WH/zGHPr8euDGNNzI9ZzEKHgbmENkGy6eBUBMPVcgQGfMBVZ
nfsPeoCq43h0JpJ9n0O90gkx9axK+VjxjW3B89r9SoN9p0/YQIV4ud6vSWcdape8
j04HUluDY4JVGQvLAHvtjwRDwvW+vz+f1Uvd+tRR9z3XMimcBpzRrVDCHRq4kQTO
wt6ZWcC4aL1sOFVfrHn4otNKaN208UJzAFKkSDQuvh0bdRAcxl4Ao78jXV7jwHID
QapyKfaom+0C5puhcKQp+uugDUNtmExXDRrj1WpVnsdALPq6qE94IzsyI4stvOgM
OzPIWGHTCMrR3cii/wadzQ==
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP15_1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
EUndqjXKzTohX0Zmt3FlcHo2Q5iCnsOjAtANZX35EDSH+gt9Ww5yZzOqUQILjzyH
8ahHpPn8eZc653IcljnVvUpfEAKnxakvU799ZY1qbxoJtR8Q/YG3v150McKouRFZ
zM2IeWhlk/9DeC6ATCFy719gmFFiaR0IoJFARMyIYGNP5Bh4qjRLJ0Onmfw7Fy21
dWwe83H5yP6xogCzS05XsdLeSSepDjMS3vv7alvS96HSHf7MOyMlwlCgxI+BRQzq
iz5LdtoB3DCnFoDexDMdVOaHu5DIRCICHFoeBJqaKli8UUsy/QoZeb0Y4hZhJqmX
90z2NaYwPe0d/O4PovvfCw==

`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 25984)
`pragma protect data_block
2YeKMRakiq+TrLyIhtZs+WZn8H5pyc946CPk0+47IqRqnp47F10ap0HFjxH4MKTV
uRfMP47EMGqsibiqRBzW6SAPvaCKQvw/WHBuqCdMX8Zdy0theyEDvoHC8N6y4E/x
uFnNgBNo8pEUfIkVlv3lZmKXiDwWvfi/WLN+ZXZAm0GqE43XNHoBX0en/BCTmyUr
dpFp7Scw1N9b1uCpG/U+qMUik0oQFSTwSDuyiyn6QAMWGqHgCWMI6tRAPGTsC2ac
AJtplFycNi0WEAJi64S4oGZfnBJdJXr1RzDWrIhcT/OQnqeNXScnJGbLBELvOqWS
EDdQVlnaEm42Aaq3FHCMflFN/4/GfRdO3NokN9+RT8cmLoqYiHnh3eoyBxyyn1Wg
YacRQM+OnxTJ116zfRgL3ii5qvp50qBq/Mm0wMMSBBtaeluMp+GNdzb3ZvW5wybp
GzCuFJy7IK+bMH8EIzZiUUXvxPtt4vf+N6kEOVRO93AXX4zV216rsRW8zax29m81
2POqYAnqX8GqJk5X15OmeY0zC66Bs4AwG9KfVDJMs6AnUgB6FKSLycjRiBdiCNT0
V21XZbeDLbxlud+LwJTY+/XeEzvkrB6ofISA01MTmbyUskk4nNQopTeoLgZboBpf
0LpGKNqA1UwxF69/cZlAodPyZJEKa1AOPuTNvsTNCLkNRMasUA+39cwmpG43H0U5
hmHGP42ExSEy7P22m6O5btyHxb3grO95/3TWcMNsKcPtHrEamfnwCyBGAxBYltly
SifiMbReFjARQeavKzpTj1E7HF6lEAlGlHpiA1ZAJecbaJx+ATOEnEfFEOalLZT/
1ywq5T7l0Qy4kfRgBGosAGnMuxGLsKPrz4rVbIBtrnv1Is6NcL0HNUAfzjFAoQ9t
csi8mMfyCCWLPN+QTD74xJcX83OciqS7H7dI2m0fFQXWp9vInsq64VEDsHO8Epx1
cnk3UekZKwBA3qXx0etX3UXEPHSz2Fh2m5uAZEnHIMmO+XIdzv/wLMwT8zRfJgFB
3I4bM8NtMZhYNNaxAkeCJJdI5CJu4RkceqQJB8rhK9ZKCsvabXYD+sU0kPc/l5Wn
dXsJxEvAv4/S0qWhi9lhZF7NtpTvTJ0MF2pk3B1RZ+RZznU0SKNQxZGnlTA0Ap9r
UvS2engALuVPr1SuC+Kw1eVhhfgJzykae69FXYFbbmhywcNBqF0TTn3mDJ3jh9Ng
clli57Twd3f49QXp3Nn8kcCSzx8LWTKSRrFIEBntnP2CZuwqwZpKDZ+T+bUMYTHD
QUM45ONjKtjmYUAvZZvkrzQqO712w1tWEGH+8ymgYMEI8449mTnd2CpLeOyTYalB
QdlyeU0cCnG+4SEPaMc8zWPkTh5L8FCZDmvEnCAbPdAhDnMuIVVSaa8CAnU/ZX9z
nIMNTxMk5pcxAlFpffWl3c39wq8HlP2ev4FT9eMhLzFq4lHvbBlty49R4wUGRfW2
YftBrm6PfUjZs94SjhIwkJK3uCr07hE6gvm7NFD7cPJbFP7kNzB8CePg8ZZeEwTx
DT6/LtOUXTw6hrlzLoWzyR646mFkUHI/QXnII2qs7Yb6L39iwP5tYQ/JWPYtWGO6
ktjrPoSUFKtImZjgdwKLD4WCv0yPd3TcriehB96iaJJXh88bgsRy4XDmN/xpVLHn
N596Ujppj7O2waoJNJN+u8Nl0NXVjMh3KiGhK8ZJYzPdrVFO4E6+RJSPN+EB0vxn
xhPsH+Wbxe+Z0IoG9eocUMlqc2q3dNH2rGW2SrBYNV1ohzNhXb4NPySnuyaYmELf
h1gHXXHfILEnBw2c0Cu59q0ZbljHeBvfOEYI2KBE/ft6jpZUAhCELf3VO3sDC6Aw
vOSlX49BWXiGosOGhUE37zSUw3np+d33Z6nZogitZiNH73MtO5AAtnM92Oho728E
JlztAF/tt7TuHRwSvCxwHWzXjb4F9UgS+C9LxO/Kp+u01uBEUaoPAF/e1LquA/Iw
9iaR5abEL/+UAC9yxsamw0JStDubshnWQ3Sw3yvLl0xB4FnFHiK81pNivOd2mwBd
HAzF5IdVwfp9Z0U/YCYCagdJx9Jtn4UPWqun2WKcJG3o65LDvg/gIs1miuUUnCDP
whv7Cahc+elBa0Pe+th2GO7K+FSBmYCkqpQS1QdhUJVoKTqya3LxSgULVifw98WF
n4s5P6+vXr1JV0MsKnaluvE+LWihTgoqizkiaPeedPhRktUDB0VS0bl8vvNM6g7a
ix6iSXA/Y3JqDx5rz1p0OLk6ud8QVL7FbiaMe4rojpXgP9bADQb0vrGaMCXCu1Kr
DTkyc/2TnON9mR20XIWQwyNMrzcjOWC4OB1YFgfvo0qIc3tF/m9n4P4D156sSbPi
BT/5IiGIcAdaaUEc2pg7l412xXnJfRvdzasTWslGkRoVphzf/soFFSVdMwn1ea8K
BOjU54joPfTzRk0S1ebrNhWnE6Cq2nFdObGr65S6ovlWY718ByuOXCAbOn8+UTCN
3Vpeu49Q3e3iMfAyq3/2+JH3MPeZpWPK3tNo7ZXXtARLhVTe2R0A/rkBf/1VCZRi
VqZUOLHdCNwBxFirYJu8Hv72BcuJfuBnn2qW43Syxt1a5CVAdWmDSFtXJvcY5AMO
gWLGSPCdv0TLP+GqIEGmP597XkXS+n8DTsodjv5IGmBs+kqhpkwqP/cPZ2bS+5mW
6qs1mMZHAjCX7WtwZ8XLDI6y5xa4C6RkJeJ0ivXsGHDwbdCyczEZhudY51RMqn0a
Q/wdP0Va78/6mKjYubS8tqjI8bun4r0zr6Q+5+SlKTRuXtdMgaGhgPzYMMqG/pYS
yMMJStKG5WZyct2f5DZWsG/gAaUGfev4tlNY8f5aXcTFInANKZdKWo+cgYMHf9pp
Pa+FSbZ++GoBs3IuIdhf8hwt3tc5CwDlrY8WAyDTkgTa411IpI+Gqt+WUA2i0dHS
/hXIlFptwrRdcar85ZBFDhO6Par5wENd3j997V0fE7VHo/Zaiia1I9aKlGnnMFcO
NrK5YtmqnRcsxXJm8t6fLAOcTgA/apM0+LUgZUqr88LTZ0ppCUXsSK+PrA8EVViV
qLl8qXy79ZbQX+C+/IdlhM1muwGpUf+oIv8XTiiL29KyXx5O/AwBDcIFGtBoSwgl
UZPFdhNbHgsphDbcoTmMX0iZc2FK3IblMehVDVwM3JUEvt1FX9wv6KlSRYKb1fDY
kMMaRiQvu5MfSGcIVIiGwQv5Jo06smtm1gRIVEGTZ1Jn7979ugIyNwX1aQQW9oml
4LIfjXzzfgLHRh8uNE14tKbvPDVInOeuANhXlnsJfGBN36lD4VokkVOcWyHztJpC
QOZxUlmsdXOmQtcF9u93vtSZpf1S94AnWWXeflerbi1+ySrXz1z37D0biuZR3Je/
t8l8zeZ0ctJzvnzMnp/MChSu1l5fjHHz7koKTSh5psuOEplgA0JsEk48VKt5MXWp
1ZZssI/M1CwdzuD3v9wPdV7DGm8hFqW4UOF7BqkbtcJApuAHP8qwJULnbDwNgPyi
WF4YzFCMPRAnD2nfrJs8Dc+s8iVVyBhZmHdnUzxMwZan21kZIK7UVi6/5c//mvQI
dT1T+XwRLB3JoiU5Q5DZ3dzo5aBEO2/WayUA5EMcSmCrEX2NEb96lHzGJmoXCENd
SwkFAemXd9o97JCWOSfieayY/t2eZLl5Rho4vPLFowEp38/c5yXppSMXsCS+IGUV
Kqy+golyKB8p7npPbbe6KYhcp5pftJsDyOJHi2ovKt82JJqP50itBrLBNFngkOes
HYFSxzVKrqirDBf2VoQr6ZvtQvqy3Dy0g2ivtdgLqnelfmCVkL1c1DE6ZricUPcP
hcD6TPcX6K90Gfu9HcNOLOZnwEY6oHnURfV/Lsm8wx4aaSiuZDr7kEee0Luyy6Ha
WQoAO4LPxrO1q80aBDenVY6q32KkqwdxgXXk+yJQiQyuv3WkSIdxVLRgFLFGO/Ey
h+goOcjhdNix71mnHRfF1czOTCpIGy+EWcEDS+m4+qpxc+8yTJaWScQfHHazcj4j
ZRaiaXkjvc5qgz07UXG7tDlKM/QEvgTM/hyLN/HgkGp9cs70SN1jn3kuCguywt1g
wYQj5xrHh2bfDEbH3BTi2ay5D//tZEukbMhH7hOuhnbJyk6NSTzLUX/26C+dsex4
9DGj6OaczYnjXyyw44tW2Q1A16VfBujYEgB715Q0keKvUv6F+XDocTtoDHJ+HZ9u
CSj6iSxtg2/ZyJ7UOHrOlH0RyHte3cYSH7qSlPtoA1Cjlzim+1muGQY5BPOzUas/
xk0g1PQgr8HOknFVn9NHyIBn00YEoXblXvgzhRbtkKonLVNgRKBYUHqWJjbz4V+L
jZdDbyeDze1Ls5T/1B3lKjSPXmwqLq7pgeqWwI6jPOL5Sy8xmtOtlX9+C39RBYcv
N0Iht/wJPI4Ealg6FQ/e2JxGOn+DQEeWtPgGCm82kwG8K2WVnjCwxkdVejptihrj
8bxywtXzMeBDRbEcnjIq4d1prBKxcLCNfIRRL2z/8ESjrjc/Mjb6snU9G6OryufC
FVGvzMoYKFMrBl5Xp4iX0O9MdikQK9v9UY3r/rd910KiBOsIvqSy9ob22djpniKM
qHK4bA1YILSC8yLGs9lHbgud5Dro5joBG26MyesWkmQepgQl7Uwesbnoa/3w8DZ4
P68qsTGbznE1KVMYOLwCcTUy2G5Yj4U2VTcUD2yZXkvBgTCDBNERMcOfMrxrse9J
L+MIxh4K0XiSK+KNI7Hg7MhFtTpeBVB/4G6/0URTaSoexiEBK4e22bdqXbWAiJBx
w/PniLBtqvtJQP9/Mktkrf7Rwby3JcewKJEkJ2v31zC5fsUqCiQUTv4oP4gMLD4p
5acD2CFPqhva3upSubxM6i/J9hogzqnUZVm1lcfkKh4qn9Awro3UIdFFNhdWFYTQ
FfCHNDu7AmsiOv9fSwIWiCZ7VVoV9PP7P3dCYpc6Ep1Tnwyy25cofsIp8TscEO0F
eYARNP9DQbwXYaGVwj2C7l2UYWrsIr0Ipf62CzQivqaHyLW0Sy4QQHbdWaW/tmwK
6ZHJtPYiksEzHnhYLk5eoQZj+Doj+VxZ49nkZQ7Rx+kkSFMnukWV/P00Krq8VYWo
t59PnlwJLNtZs2I1T0yH/ZMxzyQMcI/uZbcB4slaYLFgy68dsN4ID5Sr7NDd+WM8
J0L3tcyLF2sqOhbCYAhwuhl2xXn2Q0mLKS7V2wMOzVw1gwaHp4rvzs+jrD6Rpw44
0EZpZPbPcT8tmqmcmQocHagIwcAPSFJy/WOcqpDN2cDARDGyWvD7Evmosey9oA6x
HxsJQNNv9jWqe6NtGI0a0+vIqAf9Bj6bLgTT8M1aIXg7ta6EXQsWz932Zc2LUU5B
/koG+ysEJ825i4tW7sTRC0XpPws0db2GGoyfGJXs3lMUzyAIrd1Y2xRcoVsf51gw
8XQe7Jjp4TAyHmty4C4UPF8VWS1UBM67Wfjf2WUVlu+4GIkv9Hwqhf/ByZm6IfZR
jXHTkY+rvAcYuUZQ8i7CMede25iLoE+D9Q3qzZ8qFdz6FslXvay4Y+1YjVmzn7w+
bZ0SiaBCAZCUvOKhEcPqg6RfObbQ+Y7IIqQCoL17uD5axqPu2JevMUO9C8k1aUuC
wHGJ5nclOMG03h7X58sYsbH41dMr5ebuMqLlQh9f3PKIGvtLH9INJJn4qVDh8pte
2GUPzHenRX2RLyXbNJsvywPsVxRGxnJZhcqgTQU1FaCes7VNUPUiv8LemKqNz/Q+
4bTBnmys8jJtyqGgiW3/ng+ekdQYjkyimL/lp82yElp2jdxhKk/IrBgSD5+R20ty
Htx10t3uzjX/k0ooo7LRdEgCQ3HilWanQnvoEXD5dGHmx5CL+MKTPqdGwXi/VhvF
3hpsOPQ5kDyE2E3y18qkp90EEdW46W9WTwCR0ZWUIybAv0Sm41Z90UJunf6oMVCb
ebSSz/4LcyS1nW7noL6CrQoADBg69OcjsktmRcOMijIRTHi5xWhaXudmEubVBQYa
Z5Rsi4C/fnSLnPnTEnrrEJvNtuSddyBmhxSEq9S0SV0Jl/AUCSv3uKNm+0K3tFjq
5mCxwQWq8P9aotXyKdsqDcBbijF65dC4/4QT4s/+w+KydPZUzkjifccnNMwN6rZj
o+C5rA93QkS5VMOyl74dzIzRQo0I0n3cFQbwVOXV7BABXRkkeDFZHCaEZOWNfffK
j0UbfnN9jNrMIbSNWZP98zRFIlqFb3ctP+Pgm3lXGywwJCe4xrI7/cfIZdiDl7w5
Yr1j9ibhhejt/BbLX/Omim/kL7Rv+0ePFLxz6NVotK8cY+un/wfQDpJU6ZuKTCnK
CQu2POsGehT4LpayX8yqlGxRGLkYNv5GCMXes7nVUGso8xuh+eu6RjSPlc7DanSZ
V8VMZUGoZYzGZGWHgkZQbn+GVf33wv/Z+YHSGj/bOhKqq7AfTGWD0f62txvCyyWN
uFbSksCdEPwzXVreOqB2JdwUpf7pGywd8o0A/Apx92TKCzME82J9m+sXvr+POFKn
W6IlZzR11ejGzsBlCczRdkSJ+1Gmw68vNbceROFOSv787R23tCQ+NByAmarEfCno
/0YLfDdy8iensEA9fMUxBk3ZH9o4KMwc9U5S7EW4K+2OHLj1A1tgwB9dAG1dA8bZ
OJl7ta4BY43mLeCRSlvmNokkYX2go0zBWh9IUtMLg0VXb0+KrfcECGBA2tKPZRZq
svFJW4dW7X8M+gijArynmepy/+aU6gJnboRSggu4LvgUNTJOz93Ze8ZqYIfyJc0a
35qYudPfLAwWR+FT8RoJfgIJuLAh/oxRD6OPUfOfMZHCL1Wlga1LkOf5Glb8tpgo
Vo1Y2B9Ty1E4R44WzzBoKkkQcn3DNMGf1s+BL5TAxxM2nLnwmhfZBEBDR4KVhu1R
zFhlNsRoHZ311FrhdMaaCTMInrCReGdO9Nq3DuRw5iq4exhEmMKuNDq6CRiyk2Xn
eCZ/6C7t/OzOQxObxFHPs8ipriBzoeJQnUpIpixj3PF7PKBTWt3URIJbQGki20Rs
ZOAGYGWcjLiaoV+EjgVKEWlP54+JIV9MMFc6BwlyoXE0kEiNtuRrDSp6cd2UoNQT
lcINM9yHLNbcnKfdaSAQlHexkRJSQhv8nOZav8H/4rQJ/SGl7B9YCSiw4nrrNu9C
hiqA2USFesMTaCeSJNXxdO+uD4RoasP5eb3mPlEaZEE+CmZz9WHjhKhZn+/DeGRb
23p+B8y+NvMVqMbUa0J6BEF+j05mhsdlO6h2vWC8Sgg92DLrDDcn2dB4D26S8FLg
s8u3dz6r4KLH3fJDAAgWYZU5gM01miLPppjMlgiEQ+JhkhE4IttEdLlIc4XvdISw
SzwGqkAHKuXtOWVuwHWrLnf37EWlv0kj3R7aNFSciXmHAXwhFsCSjJuf8y5opH3h
OdS9vZLYwkNC37PyfpbCK7j/AEf/8qzYyiSdaLpNuLuP4oCMC4IQG1XH648W3xyD
nxH0Vff7Iv22HyQDFe3dIZ8ldHzyXECCBza7r3EeU/ukqL4GBPNP7VfOjXnV4TDP
53qjM60mH+rdwilWoe7+WbAJzBXbBuDEB9/RhTrVi438rVWSVvQSRUeOc6JvEBmf
ouuMBMCGS32IwfCKtH8wv3xKSDR3+RIa3y7fNlZ75fZ3w9iGFnwQ+2fEDFRWikx5
FHRCioLhHCCzqTDvLafkutfqu2G4sxbvYk2oBg+RWqQHytlEyz7uUdXObOnBR441
91Nz3Hyf1m6YDFLPckS8yUaMFqt5rIvBfJ3J2apB6uzuf/uleWu8ChCDNQ3RMmMW
RRV0YLCdevSielJvobLP3DwgY1nia4bHcsel7RBwOTSMQYPW1hnN48Fw7s3I4SHx
XkIBw7I0sqp3ggAmOx7NiAtG90+KUs76ZQ8pVl4AkmQBLF7HF7gPG/qleLyMq0ZR
APe5BzOxvFBGntH5143o3eyDmzefITAmh/p7Kak+XVf/c4piq+/YxviJof0teGL3
kPNfcp7fuVRdSfCV/DwT+IuMf7xwuCLOcDL0YC86RsAi7/ue/IsrN7qY/mgWr9ir
cPA17VZTH4gqh3ck2EM0szUcrOWeVW0EiI8/ZpnRm2ADhoEbXJnbnYqJ9BYJ3/Q0
tt9CxI4a6IH3/LnvMsDYeH3uqTXE9SGEwE4Dl5ya4WGuTIsDfSbcqeX4h2VCNs0m
5Wsp2WQUfvUEf+ZlBPRJ+agLzEzL4MnG5F9mzFDgGt5JrDIEkAYsa0m5za2hvdnC
KPdLSq70NacBfMEQ7HtSv8bFAGOIvspMJG9+UuTKeI1x7WZgM4NseHbZIWdiZcJs
e94iWSaALkRXB0yeMgy9vHnKzKm+L07WCwdv7kckzEjdAZ75/3wO41VD9QzPmD0P
Ispv7TPyYMkqtjzsKs0LEBapNjE8v4tR7ijCShMxvH1OstRemkVioCyhJ47g2iCK
9UE/Vivy/xvMW6d43ufEhhujfYSmy7eR1A/IRm87Fo4vYmgiqyFWpjbOPzLVkZqf
5dJ6NDMVqM0d8jqUcmd2HrXHkiK0K6IYqXWnP0M2rSFB63BOlDKYM9qrm/81VpKf
BEtvEjMI2mrJgVcWxU4xOcP9FgxeroBMrSkvpKAGetxH/iU2xnK1rNHBge2nzkuK
Zh8XTKoN/ItYPZTmnlfIIPwZ1LjvUUdV+JWldLQqxkwGWnfxTm8nLuGRSpBRn8Ng
IHfgwaRQw9qyNVNzowQYzPPo1n/LItKisYxbEz4U+ojc65qskT6VN1Dp4sebzeJg
jRVePcoxOA9bC65W3DVTj1Q1U0saXL2n3mm8NObwtq4tdzKrgSkVyhCGczEODFdS
JmVkU66RGs9D9QwFt3sB188S5487CNO8MjiXfJ16Dbk51OOQzkcSVklK7THjs3G8
lojUjsEFymvOWtPiLatHJmlJABJZnB1YBI701wq53mo8Hot0eMArN/+r4MQHqMIQ
Ixau1dlFv1EvTtTWQ0foJgVWdMJVjIGVycOv84d0hLHvYrTxZwW1/l44lz9nk5e6
yXbBvzdKMAMHbV8l/Sn06ZcdbP5mw808nHJ//zvnZLuw4ICNpFP0tZBiUr8RXYUy
BYApuNsvTfQoSBk/vV6DgHrQxSmru9Qm7h85LKkVWWE1ro5Bcav8w4t7usTBhJlD
qbT+7LdkEdVXjYMd4yDJ9psg3gncvplMaBalnGfLT5RCbccHcgIbpN2fLGkdvqQT
Nv9O/eRW6axkp4IGNEgGI6JRqWf0w6GBww0ubWsq2W93Js4OCqJDTOAgGI1JUiZG
1BFelJp3YCxMHM0/KuviI1k66PHl9glzvsZwTFg94JYdcDgv4hIQISM4qEQ5TUof
Gjo1J4FKM6KJtfTcNR0AlKQOHCWiNTwE5Ex11TEW7n8pyBX0AxGeuiJ1rninL4Dg
FUTP/8wA4Qks2ZTbawHRZKrm67ztv6duY3tY9oFrVaV0qs7ab+W0FOF4UYLDuFCw
HQHSEOzbnBnBt6IdZ2h9P2SE31cZzqumpnrCJmeuZIsN0AgdTkaIkGSOyAxFmikA
rYLfqsllaw2Kzwt9KRDbRduJnAcx2DHUA2jx679CzZ8L5Ub8qlXzrdN44JnghYw1
4c/Rn2c6lmtL00ybjc5DW7ETNi+QqqowGVjen/cQV4GPkUr65JwIoap6P8o7cCJc
UIeUYFzO64fax5hiS8iFmBflSkwiTnxDKnbqTj4L4JXsGFOJHk5y1cE4ToJAFJv5
IxyWDFzidT8O/B/eadb7RzIwvQLguM/rrAwuPc9JgNrxt34Sax3/JQWtLxvmzy+3
8+oEBq5yUtSAA2X2c9m7XAUuiSe5Uteyr0O1gv9EAIIi/7dEjSEBjZFe1+TwXiNz
XjKF1KhIdyXM7f/iBCkwI6AAGmFz9Mq+pg12txSNYwl6D7oE+sw8DKefCnN/J3tT
QY2iQQiAQ9NsMdrKpHCf0tA2Nia+qO3Dgh/tI9wKzYTEbdO1hBc3Qxf0uynUFTlq
YSHA8LYlik1eVlNz09XzZ4LTHCYEvr+kqkxNeSrQ6xcLHCChHW8G6tJCiqiEa+Uv
jdxShsWykM6t4A4TvZLwzZct/ofnd10HyQUOlOkKm4YQSHph3k+4dPepqU8ReEBb
UBxTjR45R2e1KhYUsF0MtEmvRVNqTXRR4e6t61lc96DEZJBWKpw2XjUSiRIDXcJ7
AwLosn2/VogJTa9FDCp1ornPUVnTDTUyK5D9AtMk4qxoCPCJvU8n6BI9FRvu7VOB
T2ckBtDLwn0ggVpM0Y3M0EyH603BznGOccs0urGR1xPmZTfT/LW6QcA/N4wCFDMn
wdAKRUeUmGlgtRKmnX9mVPRNcduqaJjDR4tXXy2IC0YUQz8kyEjAuSz/AUASbYMZ
Yun2ghwrmhOu8D86WcTWyojVKf0RRxjOSX8nk5tEtBeYuj8h07e90LTRJZyjHZU+
+YkqdRDzF+B4O1QZryPd0B4oBs4JN3c1fq0I+//jYW25r6o/KnmIjtL9hxgixBrH
/LidqcKs+ZlhMypxe4S7r4gIyL1zFeVKk1R4rBld5QJciPLcvmNkuIOYHreyX5Ht
TQJ9EHPPXgjTcJM5kYAO3ErkQ/rT5GNW0J/Umwva41gSqSU7ZokuEYPwcYJ8pHLO
4ySwBYkB2WlGeD/zhVWlV8iGYnqrbpMmaX/jTfUXmqL+siCkdrtEx/2aODLE/BNT
2D+gmq4Jy8ju4DHJybCljD1TL2Ng7JN7ac6fjoJ98ImG7Earb+h3noWATLMSyKjv
4mBIN4MIrdbCPp2aFVW36fqmGSgTDTj1iNETg7sLmT0ttfMm400Vli+QIqvbw7+F
SJgzZkqKMOQ5R9TkfoXtoZrO2CDTqyy8Fs2/rDCK9CV1jzAVCgH9Cu+Rz1CrXjKQ
tjMASsuZXhRo0crDnMUF+fZ9msWyjQgTiJX3hjHXlmdv0ZpjrL1NIXPPVBMDU6wz
A+Q//cTFz7I+ZAVPMUKjyvnNzNdf1hh3kZXZVEpbSPFOW28pVJlWc16vnTFfevhm
FKX/vvnXnfrWYmjfxw0Y+Ca72WBi2o1jCf18NEzva0wnxqzQj4TLIDyRQKt4ni8A
5EBvbpBvNIEa8OfABgmlPbQzBZPHk3n4Cbv5QMOFJfWj9sVw66rH/zaDkMF4szbM
KS9FbGYlOvMwstpTSOeU+gXH8AJpK8+Yi/BQ1nDkLHPP0jgc4rQ4FHJOI/HO8k/W
U1DYi56mQq+UEHuOUN3ZkF4+KLqnBzOK2PmclYz/eM1AhJvQMM8o8c/eWOess7gt
r7kBhuHkoCcQ2w+ngbsPK9Ql2BBzSDpmnb5YPuau+DKQvypZGVwI+ToqgHuL/+5N
3z+oJNutrMKF33ur/ZvMndvACsqerfJuHAF3m/cEg+/Uh4NZRkfH9Yc3PsuRv4XR
0gGf9TBWRIeypXxl8sSbvDJFu+NISoKWmBn/vKGsCf6dklgMPG/y7oSxZ18nNdaW
OOZzTUTQPq+OCdEZYqBVuAWQcc231xjd/4nB9JdRGpJ0adY8sOk9n69Wnhz4oB2B
DlRolge1Gn7BEVROaIBRV+aTZbTUvQm93Hjzf6eq++hBjPcAiDIcyO6Pu7U1w9uZ
LUW5WuKWwu48iCDpLZGZyaPH89QmrFNmV6ywuGY816j9krYdnZ6i4b8XA/iWGt28
0gz9TfyP1scN1KkK7aymE2T1aXJT4DCIm+aMQ5vflp8bkqQNGJ9kW7QBR/9QPEkm
XtCmA9bSvoz35tnhtamFAB3HUMBrIoz044UoYuOYHeTKlYz82siecQIBDIuRncZh
rTFgXZjCRBhsjEHdVYT8ZzCU8o1YAr5ITVcrBOe3bMDbPWScY2HBUrdliL8TtTwe
LiVeAcjriC0FS8LPB1jiPvEi4pw2Kk0CVau+D2A4O4l250sB2C67JBpgmPiQzXkV
oJF76rsGdZp9buquYgaHHiJv72AEOqAR29SkEaFiWUUy5OOgQOGhJql67I0gXqUe
MP9wGh7CY2SJX55xIloeBwTPvsRy7xFItfCBbk5zyXkryeB48Lk8SfVAUg1ivjde
9Myqz3gMdGSFJHBwOF81bCSEV05yBu0gXUelhuo8E95r4AiJDbGCgKwKW+ExXban
/v6gpZKTIlEz4f0xz9ttEo1U/5Ec/+qv1NkgrbSh1DbYzBIYdXcCdKF/MrA5gPFU
6IrHkBhIVXgMAMiXGUQaSXwHdYx+tBi9Fib6VoPuahf0GTMaDUGv4yKdEF7v/cVx
cE2wFcnecqjxQd2iHkVfCxXRP4/rvHEa4FE83BRXwCsLsdHCW1neJgLwM87DMsmx
6z4mqRSm3TIbqKlYI5sYW2WgZW89hY9gtvgpSY3kHtAMRR3Z+aJVN0WHkJX+njnN
ZW/Tj5FOZKwW+KK88q25Miai6fuWTTQ18QPGB/xrWNbarhq9UiAhLugTRi3Ck5xP
mJiGI/J3n/WCBnJNK4KpplbOuP3jKu1zmL8cMWRQvgdzQFCA4BZ2iEYMDksgBFe+
BrvliuyfSr0pt1W3nz/tFYByMOFJQasgvEiq/YRPNd8OBZ/0YqYPpJ32ef2MvPW1
biwzD0dk69Poxn2CW2BDZ+nKLXecfqyasT/uBkTuiyBzs8DWHsiiAGNx2lfoBNHP
YoznpGubd7H9JGjPaTvBVQSxvYVICibmgjKv3+aw28PyE89l87mA2vmeazJ0Rf2c
KxZXhTieBbnzdmS5TwbgVCf90PDUb7WgaPgYPvP6WWfci2gJmkB8aSiJj2DR0J8s
CnioD9JTfff5mjVLsXNyQJIpGSb9RA7FS98uPyh5lFWucdVkhkAGc+iTadaom+N5
LKJCZluOad2g8f1ktTznLsNhv4oekxm+jYEBaB7ia9ikYHeLMW+UmFQS3bQ9XYEc
q16bMzczOZF3GdQJPVNSvTpTCoNLpCfjzO6K4x3NdvRy2ewAsRXk/c6fTNaWV3YO
xfkC2PKhrpySAOzsgZ3HpyEjW9JuneNdMLzS6Vq/AzFYAEy+ke35KXZTGSLjd9KF
2Rj9rRwwXDOO7a7hkMCYsHdqaDasEKQsNX6nckEgaDzTOA1SHZWTvqwXeVjSfWlw
YPTh/bPL7UAmP/mClFrinZiqeujgK2tmBKGBYHazpwy1t+MXym1ZWJ32abkR+k38
GVDxoK/vozNqrUfv0D9o56GEqMKHv0deohaX5FsuH6QzcGWSrOBpxqtQ31BJCUFe
UEQb/0t3WylbhGv4nt8AiLPN+MN3rT+5V9/CMQ7RoF1ub7RoWGnG9r5NBPzaSAYJ
quNWlPp93I2hO7jjvLAgAqkfzlAGuVsVW1dY6UMfOPKW7Knyap2lTEN/vQGYcau0
4P+eIvWub1RL1u6eT+2n8Yh9TxGqfqTLh55fudqTYnJY/M51MIsgVmrUUrHUs3He
7QKwuIuDKIkayypQMuAagVgyuq8KWnKdlk7nKC5SWLIQzr1qT7wvek8ZXwrmlDJM
jZJiuz1cqhV6W+MzJUjSiKq0MrQ6J9KSbhzeYpYAWH1BpwXvegSKu/1Ts6/GbjTl
3y1P9qLHfU8v8QYdgugl4yyxqEEJO7P1vQJNcU0IJj1Rp+9ZU0I8PLHkSsCXWpgH
GEZzTGbYKb2my1wgYflHc7u4Zezn34ehz8JGInie2u3bdAM5dJKGYa/apUX4aEtK
OytrIhXWjivZOQU9XHtAgfrowDVADz59CqyKtRpRsDoaoChkaQqGIsKGU59plmNb
ZLtCrQwUjjJ1Nwy6v30rIxacShUFNXrC0leGNJKxE35ACoiWdhWEERRGwlHDt8Nx
CdKU7pZ9V4/z5t4oyC8uNTZZ0buNSyKr5zBttvTkkpYElDgx2zVjxS3R89+JAHm8
1mD2sMbIH/uHm9ViXPanr9cnGXM9/5WMW/EJtzo/OBGcgUxPuzTFUpuccgCIbYR3
hVO61GJXYZ0EGNZXLsfeoxL8cYeUPV3i8VhwjhXKoTKchWniw6yTlOCq94E2LBwR
+WuQvxQVw0/fvxJ52nPNVIACXsJj9s27ptUoZEyhxdgrjOwTYU0ND3pt0xT9F99f
0WMKzsOSfVBWt2YpuubFXzD9dHH1W56PMGmUDdbjt2pPd5mjLYFSlVMjzvLG4I0A
A0rXIbPtCC22Jwz3DLFMAPurfIVsalI9fMhy+mxp6wG/rSs/fEmhtmTlAdRErYFS
bhoz/v3oLwe78G35Ghe3OvVTLbAnpEBV0xWgLC9C3JwQPrtAGFZGQJ3QrJFk/nxH
X8hvUSKrGBHxMqafwfcANuagPe8DgdCmHHeL6OKTiI8d+P4iXitKJfdZSnVrzd/R
ROnAqvAbOEuWrjpIyXqnnfeUe5Nv7fBF5JzROATZt0Zhs8Wa/NKFRH1Q9z/0i2zf
fE9QIRtCNxFe4bA+0lDloY41a/doq6AnBSTPpBgsn1hq381Rl3DzwPHiet6zBqDR
3lyWAkz7KkiwfLOyDBh4eTwnndfxXBvgt0XdBiOB6GXizfc0St0yP5Xsz2/4JC+n
AB2rjBsABQ/pbMlrG9uvB9nM3y0vwK7qvdkREYTaN7ccvBuj5a8IdjfZ5KRcc/Bm
XBdL4UVyuyJhbxXE9Bkhzh556jVYipU69G3E1ruDXIeXXHZbl1x+tHD+DKbWxpIo
cFknWmhrI5uZKF+ARnh/zuGKT2OFevK+b26jmMjB1Nbav70DEJ/M4Mqo+1EBGCYh
npGX6kcvLpggFlzNhBUHnngIk3rK226zLFp+ClbcF6LbU2J57tusrhRbZNTSvkbX
ifi0eHDLdt/R2mAgjLeucZaTUFMsqANLBpervsGYQdx3d5oGmikxCkTGXXyT8Cl/
Sv5Agx7V8ED/nQ7ic3hZ0ayzUgCL5xTy6+zRIJCM7aqL0pi7AM1AKBpne4lT/Lzm
FU+C23zQ00qvREg0j+3n6qcCCtQ8NhsZZa6H3kSbDcIybp5oXU/vDMs4kKuxJFUk
GdM+cf0sufhS7iKPKkt2tvFYegIB4U60IapraLtuak/gpF/dnU7U7dPpLczGoEmH
0tbEfu7DHDZv2qlMefn0jZDukOCsYxTGmGoW70GCpOel+4ltAgxpALaMuo+e1+Q5
TXjxvHmQcUvNoEha+tZFXhYRGC40kdeEFSlkzLrjCiaRMR/Nv0QiTJ3FZN1TquQh
Bvw3gmCpqCuSF05kSRnAppGCCjfGrMdVRqfHrXUN7C3aBeC9htuuU92OPZdQsPhg
k5Dc2QzkKkvO0r1U9qR3e91Fg+w8Fg52rpU155f5/bO1/woQYxu5eWyOX6Rw+uAF
eOpy19/C8LH22ShfTHu7CrC8T++F74HiD2L+lHL2NltqdGIXb45IdcsvZnzSY0QL
0iabJi68lEnjwYl9g5unxPb68dJOhfUv3lw9kRRo8WQY0JkN+QfT0dFLJ8BveT9Q
+9psXJr9mTfs1XSDZnBx0T6Vhn7hn810scu4KQIuWiTJNYjkzQRHs9uxI7adArZS
h4XDQLYWK3KUauU8GGJIK7UmD6zQ4kuEVZFabCZmlT9lo2uDp8IfPiefrWZ4Bmfg
tkRNixWEqmWuOBsXw5LqWd6rdUHbfLVQVYOyUXktW4nTM7dit8IotyGDtoAPgR3s
0vx65MhPDRgaFJHH3QiO6/guK6g0+IGF6pg6klMdaQnqWmRfMSrTc6LGbbI0tyJ8
1HA7bhfNqzNLpNKfAgCDVq/S5mOXFzqN6ZpgTHGiiUrQW569aKC7xzW62QVlKOdv
jZkg9Z6Ktc3vmVJsh3n6Jk+L8IzVO1+oAZVzYJ8SqRS6+Gr4Kqw1WBFYc45eEK/0
fBG6VJOByu4bP7JGw5PGbX7dNaoZed2JzcHdv32Cgk00W72NxgVZrxpV+UnapnPx
de68+cVuRbFYcEd18sQfAG0hmiTxDHtBhDkkJnWHpd1hIchDK7S1jVa+wbHY/wYo
eHbwtmpFa9bdW7cIPvZF1ag2g3JPtRAyo0u2/hNMtJOTFvyTuMyCO2O7MWZW/uWx
AmqRHbLXRY8Gx0e061eJUhtDUXapM5R1HY3/xaIqO1dIYUV2xlTYny91fXaewHJn
WbivDgYAj93fWvS9Zh6Mv9m+DQ4I1zs96MmRblbX5eVb7jVVu+rrikpXo7BLF671
/wu9zLy0sXbaYS51Yn0b+GCFumkm0BXEZ72e0/KJifgV58MW+QhJ42C4WkeMLRKA
aTEFwQA3uPjTPTxhM1d/eZLkMwGC/PZIBT1DsuUbLQiqPDUIbiGkQjHGo1dH/SKQ
qPybHpwz6oqPHl3QHXEoGz04286jJVTsTu8ppMuEj4d87zk9T2owG/9VfOuXomWt
rfZDf5OfnRv4xdURXlwLAt9X+yvexFTuadhOiKqygZ8o4Nw0wASGJ/DCkkXYM0yy
8d0+mho8+n81syhm4BgC2ERvEpqEnC0qZQbYWgJbwIci9mt0Mc14in8uXuiueQEM
EjhY2CSL/hgEsUvNO5pt8ED9Q1w9vpzjh8I0VhUCIp9NRzfxUKcSRO4e2zKH0mOo
q9ndiGjzr9gAmD3m1Ef2luudc/a1xiJH/msArpZRQNxmrX5C+QY9nmppD6VTp0vn
Obq1dBRYTdIwRQax/WrupyiRx5fLAYWllXYTX8yp20h4yM0869i+qVo8eEWg6Ro7
z6KnViD7d+wi/pmLJUuBK61J2P1iRKQC1QWsz/zK7ZDS4WNGF+2DThWvY9rJ2YIC
/eCZE7tsiE/yQz7wrlqWvibOW7zQIm7DJJW5uASLjRyUlsZ3Hs4gIsiTKu9B1JEM
NuW5uakV73XA1cH0sxgPp//iaxpPvZ8AgEHmLDtyO8ubr4iWloyAk9KuqG5IEgI8
gGKkhMD5MLtbOMxa5PGl5NL8CXdiV/bqY1muzrK+2IgU+m6I1wJxdbdhu7ex3l9D
Al3J8EVmaSZ8u8nqK8ltC5MuIFya9S0S4WtYHfQ14VIbYej7kHOP1RdPlDiphCc0
uutMK3w5Dq3zzI3Zs4qBwNLkq6yA5EsK8oZoDg9M06hq6/7MJb0ch+P0CZb23GSQ
U9GalT1lDEm4cuLErz9wOmN2TTgdS2kOx5I4jGsdyZJlPSoMFYaHt1oSSdgURu17
THHhvDjxpNxt0o8egxm2IaloHSWnIUU06QAz13lREee7Xza2CrDHd0wQcE7olXQr
AsTRh5HA7t5zAO58JVENDbPcxB7LdMOfjN3O1wD8jOuiRsZxBQzyfpWfcrNqWrq7
f2PVoyn/IFcLfp1qc9oAo3Q8A9hsZ/IePFKSdYeKf9TkSRNDwBJ/7AOHZEy2ykyY
2rapDuzEX/VoZSmTzi9+Atk1MEB+QrV2qm8La6Pi0pdmJaoV+7x1OJNIyn+XX0S7
GO9s1z10BKRq93hAitxqqRm+AHLfAVJBM8S9SvFuPWVMPGE7BJlkgBPm4l2O4Ykl
jt7jUobDHp1edVyot4yrJnLBGWi/WXlV4BwQt77ojZ7nAfmctK36L6kOqOI5okPf
zXVS/zlQnvRGsD3GbGxNEFOzKP9FDsUKV+hvAHAUwqrsMnKqBiVrkrvVb8lmI+CN
9SW1bmopot2jINYIjWSo8suNQj2xDxtu8f5aSlJlOoUN7lLNADEVeSrliDpxRBmJ
1kmvuuc/ZfOzeVKZ7OZUa8VTmvP2rw0nsSRIBdL1G4RaK/E6MxP+vUVcVpo/PwEY
ZHDlaKO0uyt2iuh4gKe5xny6rPi41g6ggQHGHGTqD8r/MPwebGNAgdv8BMvxCxu3
PF1jfxVoEFOGC4mHtczepCKGMrssh+62EQd4Ty+z750hqENd7EztlZdwF2u1VaWf
wNmQE7PV+NPogzkvoxsLwQXuXIDVjABPprprzTKLfKEv4j8VIWwp3q2gHJpiqeQw
3sAU+I4zMpJQH4i64oRq9SK/Omc50KlvQSjqDGUViC8HeBFaDZJIT5YLZ6NK3Tn0
66kEu28US4Y77KRa5xiV90pDhajrtRVRDFKnrxR2KRcrSfDeEnecwcBs5x1/TB7X
o5W7bUdC3tKLAWGbhv6gCzSMZCIskX8RaKfWo+7whias+0z62lMurYOqXlnoRKjf
0vyhOhUSsrpwu1/eSI/0b5NlIC5/eQHlw4qKEB1DG/LqNI+aeKTRPtjQ7iQrvKJN
p3hWYrAnJ68WC+w8fJurx+U6Vff7z3FxZR9vH/5Y5R8YiQiJgrjrUkSk111PPf3J
k1wqVA69Ks0zRjLVxRK/dIQYzTcrksm1ojRAIrXVjucDzzzrjjGltJC25H/UL3RZ
PP6TYJX8Dkj2S2XNRQEbapxhOPARdCkRBmMHLcIQ2VrQqb+DH6yAnoez64FCO79H
wmXnqH8+Tga3a6qI02QxbyzrWJ7cSL4Chcr4aP+QdTuS5xSwNvdnoOxAPTE4B7rd
1q0cn02Wo1Rh5D5nqadPJKVKVr+CoVuc3RzdODV0FEOyWj4HrBWklV+mc6Uw/Y0j
UcMUscXAcp+iSvoHpMx3wKsuef8GarA5fROFQZLlYyP8fPefpWzogBPI+Q3R8QnO
Qtuv+C6DVuJ4TixAD+7N3wWY68N0GfWFWMbP6ufEk/S6OnijQy6AP+hIVQW18Fmm
EwCT4nUuYLWhurbUi/CgytsMPBCI7j3SsH3K92WTfjip6QvLo4203ADfU1iKQ9x7
sUUksQkLsHixwPQBEAM860C97V9m9oM+HksOFIbrH3Pnwk4oz3k6GROcTHfoh/Cn
EebXq1OWG9yKIzmUutXmRXhMgoPZAN4MlT6PyEIoLADbdiQlw23i/KYXtZw3kmCb
em3Q2vOd2bXTYLNn/Hnn7v00cKkLmzjaaqSLivBktkuy+QHrOjq+y/KnEbceLTLS
NZDbJZOhDdtEhM2gy42BZyI0W2iYW8OXbEtRzMxdCMl9TMuYTb7yYnThh5rgQ7uX
Bdvgex8HooNvry9ymyhrp69cc4LH6Mo05bm24OdxQgUy1Dvs4XZXsEUP2Ad7z70T
mHIYSf9e39r0u5IwZ4tESedHa3lSxqcRPODl9VDvDhLSFDKyhPHy8HCH0fCtizFO
IYEISXsl6B3mUl2u2/xZP4WZc4siN/O5pfQSpmdcdND4WGcg4yANlQCbprESL6WW
RPYOUKCjIl60QjtoZz/N/emeCPcqw0DWVOlxDYYi0yKoa8YHyJNwvBzlq0aOvG1Q
zoqmAtRpwRd5fGG3RFUwlx30pogFW4IXNhdvypJzxWY20UbjSonc9Mpx05XHoeTO
uq5lwluEDZvoabs8D2WSuwQcm2vdJdflfBbR77Q7AylnvNyPd6TV5Bd5TqdzPcQM
6DRy55nNGOQEqjbFQBr2f3FGLyjyQGrIDaWQCoj+B+s7g2PTOh0YFehzByqMjGgj
oUqNQg4rK8uqA1NAXVqOoCd4U/TwqUMltXFTpNBFZF8gRlZ6e6y3QOKKyGwy/Icg
2xxLMtE8WeVc2XnOdbweHP+b7gfIvUYE45zQvMW0B+dVOyCtICqH2Yw6V0425eom
Dkt1NeCnQobHzdNISSvjw5tE9Fb1ruOvpg6QdGC2I6dvLJ5AEWHM6F46DdsdhLr0
gsXkTxMoPkOWojPIHt12hLiHMh1hyIXlk3ySBmHt3KiF8VGDFQNcopasC2MvRfL0
lnke2zeuvf6wJ01DLWDhyVeCaMkBJMhwgDQBJtOu5KRE66or8puSLfLxwTdt3u2a
Eq7AM55WlwBx+AvALX6/cEo1/So4B1I0+i5GpdX7594yZ1hJ6D8+C/dOHjKCnUku
Sif25vjuItJ9zyAa981769rrbYrUBgeUpa88pv0oH8c5w6irRZQftcubYB2DcXx/
Z5JF3u5Sj+BwHifEN+/q8buSnpfd2GO2FxAzs9k4c82WYFXFXWqXGoNpAab1Ri5P
TlJDgkQvegbBATzD75qZFNE/IBjEGiLOiw+PjMhon7DD3E7bw88xFXl1vYFweAn2
XDw0MilyBLbBfQR0Behmeg3TBavbCbl/ptrfok/rwO1rOT3VAKKSwiuDGfgqQMcw
fsFwY5VUAx5tNbl2sMLGYV3EQ6w5e0wPVOzzyVFbb0ahvIbIEIbxzDOGQDuruUmZ
6bu8j3guZmH3+ZZ3waBvMJvp7rTRoHVGr0HWUaEjtBccz15/pg5EVBuGybML6Uh8
mEl6X9B6hRq7iaKC1kWz9HcaChB1YDRjIeB1VxbnDtcB9pwgmS303FHUKB9eKK4B
iXLZe6J70hnZbUUHZqJEXm2q5t/Ifejxwvxim+dM3pB0A+w1clVtX57jE/S35ALS
DE3yWkBrbXtp802zUslsnI5WrYHGQN7QLuTjK6AxYw7+pWlYBmV2rSlgalQdtG97
WuGSaTzT7TYUHUxRC1qdp820xgrXNhp5luN9EexLIF3f3LSFpt/TLyQ1EmmTRdHM
YoWBZiK38XIHVzV9tFzvjqXO3m78hsrAoxF0OF1qNK0M6rZqc5jbS3tWukzT874M
AnMKM2ntmzxwhuqpgLwEOBnsvuPfBVY6DE/AezFm35oDXGBqIcOX4RpRQxOx7ICX
nfsOLtWGkOPmgyPfUiziTJszPDqJzbkS5lshsk7Qq93PfEktkqy5VDQbkMj57idZ
zQM1j/T65zojx5mtb34OX5SR+dG4rUYPieB5qaYlA93ksk7EyfaAVii4g9gJGId2
fxxEiQ7TffNKzcEZPCrEQ0AqdTIGSX6jGIQeG/DV8eKkfzuNxcD75iQ5asxWSuB+
A9+DobZo1I7gNejz6kx1Tnq/R1TYFhSVnJ5eOkvgpZ7eg0rDVnZ2rwa8d/IuOiXT
vohb0uyH2djLx5w8Q3I0CrsKfjft8xdJby+X4xO7UDuln/hfW5wg4yNrPZZp3V8V
ztVyq1he7j1l2OiuQQdANRd2ctGuNVFZWIgPVfWNlZEsUqYMNgnDvIWK3eY78fxS
aSZUXVRhjRnnqUBYAE9QH3Tl7yhtsxen9IUbVPQEyH0qcaVkLRzRSqKfSE3dL0fW
VhhuMzC++v4ORrzL9b/pqyPqPJaEkm1sXuZTZsCfDY5YE144G8wnFdoTml2zXBaT
YKLbbg4ijU4Gdx8CroVnInPFowmEApcxwqCh2poMgUm/F4woiiJjg3Va/e8U/YQQ
zpT78rChmvZYYU/A4m3mNFmQLR10YGM/O8A/z1NJlpI5nwlQhs7aWc4yMoSZbAIQ
wnTOB1goeR64LX6xkPzdEU6UeCIjSBwKMSN254oysdyhpX9EqO+4+Qh1zq8fdf5p
DqeCqPwV5nWGsTQoW0yY0/Id1RS3RblnEA3qf2GQa5EGprtT1Er7qK9ht+YuR6gO
4WaVxZ5NJADyM2qEl0ttXpBaqTB8fW0l+BHEnGpyol4kk96zrD0EWv3wXWdBzglT
XNtKsHZthieqxZar9fB59zPrd5STN3QUWoo+MHnUpdVGKso+9Og5U+0z/4gG2rMd
OHDFm0j3vHFPpKcyyC/WuK3zLsuwaprGwW2gAvzyy8aJE5o3X8SRk2K6JttQVl6g
oJdW9nFAYsULSaFdDj5FJsCmwTQhN1xlAkttSTwAYIxcIJthGcxtPaxdRCeuD8e9
kdrI9EVJUt+0Ih6pBVM/BzaPdLEJhUQtkaZWy1PMUsJJL5mJhMVH9NHPnaVupTkq
0/4ioM4FqzGR2lO2uCOh6cv3yd6woTrs+V+XG6I3cRifKJDizNqYerieK5xhS2uL
6zSXCXEKZ3jkfUxcLOe2IZ4ifYS5payLtTkzQxUOkIE6pIIuF9bFIz/YC9G3TAWp
p9J/k64PBR50ABDN0bOaKtkDJqYyuTr4UHz6Ur5QkJX0tunXMhH6CD7IwsBb6eVk
R8tXCHOVAbEajuMRWoGYl5w89DqFNldCqEedDVPeqcrd6lBuv8zaPiHSrUSLycMj
3X+3MRcT+AZa3NgX1gaZHhNUQEr/T5oSfhVLd9w7Ci05KuiZERCEMtoZ3X6oV2tn
77O241xx+hp9xHlGBKhEENcf1q/coVfqGYPchg6YWhQT0KeDzD8UDUJ3dZjhv59B
2GuXad1wNJonFoMFLg/NsaCfbEoMXi4ctIkPs4poowRwMt2UNm6cDDxE2AwFU7je
lLBLeXLAxNIUC3q9PZ6RQZu45ux04BoHgUFZSSBW74FypVpQB7ZPm2zmtpprjw+W
tSilAPYaQTE+PV9tbpynLYC5sQNYSfEoSiEUhEumv2hRnVe0IM6TdvqfP3soIaeg
L56ZxCQwXeiCNyoTWv+ATGLhU0e7/Wz7+szhMkWMZP7XpG54dfPkVWju6fOGKDrZ
cik1Q9Bl1VU1xYiqKmrAERjRgSy1QJkqJD62Kb1SI+GdpKZNp5lFx7kJL0Ddn65p
ComSdukyJHzUEgGvkYMAOUrwGaNSr6u0sk7AIo6WNTHm+Bj2PTLPbqpfOvN3+A+Z
OzZeJwJKaU9VjvQSi71prP4XRaPj8yQCMBa9irmpiSUWEYv/n5VUaxQxnid8ik4z
tEGeVzAn3Bo8im+BK0Q4uKvECkOZS4C6CJYj03SpCmzaE/88rEdyoGs/q6tgCt+v
yVlqBokVqcjBLRwM+Z1d6SI66C8K6hH6I6RldwwfuTgffDR6+Cw+iwY9nrHMlyJU
AYVWcCSiEbAS9Te/jzsHZgYuYhXq7t6OLY0E3g6tEAYrt/xXnCFnBcZu8HQs75lG
x1qa8E8FH++fNvutPaJMCA41bf5F1rWIULmEngs0moLdZeRJZQuvPKp3NMAXBJyK
8QHgwAGLYJxfgoNdQu83vdiVvkwCh4LfFqVpDG4SNRaLddSTvyDGu/1z6DnwyyIt
m9NsK8iZp4lBSzI80cTq5d53OSEv50++v3kNHIctYNHJoztTO1eNobxrTkU2uhsP
LTtyQwKel2dBWd3pfYTkXOG5gnrs+lqzJrtSp8RDRKQyebHXweW5LgkwhOWYP8N4
WUsgO5dWnxTqQPwTJZtkSRFAjOaySUL6dkWWS9xy8bfBRKKLm09Z2aRmVtwAIUkV
oEywQA73BHByTuIXGnMrlPra0kZ0DoXLCJEIkNguxbiQ0bzsKzEufPDuCsfpP+qK
Gzqq6c0g7uYKepYUE+b6V7hBgsKF7m5F8u3P5xioVVYGUZCLA4xOCv9MYb0wSgyN
z2F22b0ufamzkKIXD98bZfzuW86HAEmfX46RmFjaXTnzcgElAH5+zZ7VviA5N/EJ
/UnVqnwNcu2hb0n1tSHK1XGsZNJM1juhOixhsm0t0rUzvj3o5j9amj6Y0HE7aoxV
mzw2QI+MV1zzNNHXEZJpiLBqjA6tcjX7GIrAGXMzR5lkZPJOJcs/WFYRdusKVcur
ELFMwuJZSR8TyekptJ66+zSbQlBZC2M8/vCxx7avAzeuNTMWwo0voisIF+x8L82Y
P2ZPzFTCSWnGfqIleV5NTCXYbyl6sMvqOJiwrz7/67jNWR8XthhtngzPCooKBPD2
oIe2FMocDEkqsj7vEL1tupGDTHSmir8IvHjJx8OHW0BlFzBqmp3s+39u1Vvc6P9g
z+IOCBTsLGf+ETmT6TsUsZMOo9tIFFMw1xwbK/7rIjXrYbdP5NPtmMcVHzw8kQJQ
/10lqOb3EXqFZ4Hh/vDurbPBeMET0+kKnTCWPGsA+vccaStEXzxlOAc00XkNtuE7
LZ0Yhg+PYht5FRVuQQ+gn7yTo3qcwlF2AJ1noreFrPkFKFLzTvNAssoAFdXq3qSI
Oh14MCAGbZxajtB1qdIiXJKKjGaIYC+lv8qNMgxEZZmjjddBdIacqmv/dkxPEjtP
y0qJwYDwTzB9XrILWR6YAWbWxQQhgBEAkfHJExWlPz1PInDNARbyySaoiJ01GKbx
x/EytsDsQ2HL3xrtnzyEfzS6vzah3+CxirbHW1BgN93Qaio+l0L+xCKb86HZ6XEt
9uvkNjZ1dydzOGsa2E3N8bF1VszUbP08x9EBRxkYJjZ3Ub5s5huY10NDPxydgZl7
osiay3ZxIEuaxt8ozfe123pcxebgdxW+oDs/C1sWTmOT8SE7C6BHYRfvJEO3u1Zw
HqFlXpWqfDhm5dfkn016/5a9ASCQB3Rl1KJitqAsJm7NjEJGw7Ndry7XwvmDtZFR
Sfj+783zHwDqz/ia0ZvsEAT0m2Ilwn+sWvETFk8NLD84BniAdkguIZEFKvuRN7dc
KwMUuzvFRKUd74jg5fmHeIG8/F1vljQnKdZk8+yT46uuL4SBHGma2R3OybiADmX1
TMpzsI3aM13AgIL053b+EUcZeEhAUT8NpGQYup0NP1zUWTPdfjf1AtDhHlNj5W4x
5ZiD+pKPe8GZTfPtDmhlAmRmyZKCD8oUNO+ksnBWnagvFvVDFtvqZ0mgvoFgdQY7
xEFAtsnQZpq2iv+a6VdAvpcHcwDVh0zD46KREdNeqnJO4uju9Jz2hEw6RwoNLm//
KlTjE0MgCDZonH540CC72tHH40xmPTmgOGYlOcYTnxxNLXfnNNV4Ngbuns/xFPio
OOPqvgPsB5TK8jszBUC0iJqk7H3V4/9TIGiI//i/2RrOX6dNCkccdsaYdcvdUZ3i
injPQ/uGapaabjAGdodswPTJdBK2QvT1AWNlLA/8Y/Tkz+gS8Iiye5JOnJKEmp9R
ZCC4oYRxdlmlLINwSeyZK/AtNcGzjCQz5wSnvh9LvCdgXexhp0PZIbZzxD0tGPjL
0/DZQhKAkxJ8igOjH0ia1hk/8v/pUl4EYtWLj8wEfxnNddSVIeHD4R1kxpApdgBY
RdUw7EBfBXHPE4ModKGkBTPp2jUusVSuBLX1ogBVxUljC4CGe8zMAfw2dQxRvz9K
Mt7jEohkNDCEN0oDaG2IW1kaXO7fnSJcjAhMWlTL6G9/ZbzYJqTCTmMqLJE9hEjF
A4J71ty1gFoScYcjx6xpD1E1+7DbiK7SCSX3s2TyvWRuY3phCU7S+dSKz9GuNYoi
9Xh0Ye2UVz4R52F7M91auk8/n8D4atjudySWHLTk6sQa/KzLHzdtx+HBLqcK1FXE
2MIhYcSrqQ/0tCMXfUSXo+9wsrDV6nADtqWyAbqU6yE9I8Ti0CF4xWxwZKgvQC7E
iftT18cvuepIZII3QWZ4qt7E5VJjqVRe8+XoYBFXAAndUfUdWzSm9gZtI6R65EDT
qlpb/rsnPIgwM6MymCpsss5TJEP0YKS3HBmHJLyRePhcrMwYH7xVqQ9CMsobWpV8
G1abBHBjXn8p2GrI+jXLg4/HCx0+ag4+sX7BtJf1pqwHzBNQc9iJzz6eB6frHqlr
fN7lzoWvnAgqa3uHLgcVKwFruP50f9IiG652tETO6a+uxUHtl7XH66qtMTt+NM39
ZugHIwciNGVo/bsjqyPMaQGJOFZgpVfr2aIGV1W92ZJ7ym+cG+q1wTkRTrB7y1ZR
uBKiAXd4oHzOhma+0K2xDHpn44Lg2jOBP+gFP+FsFCNRCh+TFmr/rxINv/Jh4Yt+
kEIBTNFZ9AQ+lc5Pu2NuxOl2NwawmBqOiVNXkEgAmBiUIYQQVC0F+r/g6JtFsSWm
2YcS9/y4aZVepw+YR0LXlRiFBNn+mYAESFRKDOyLP6sVW/cKBPhN5wr3MreAyoqL
q/87HTV2dZ0hgP2lrsdXKVukI9yOLEHUboc1wlE+y9V8HCbSKvSnTTlecD4qd4B2
1XcSWWIhEs7yapAsqp8gvvAx1qsCf63Kb3GQQgtaeHltQsD1cCGxYsPraQufZRVN
d5LvjvnUWUYOuNUgww5GP7B8zL2yA8tINZzW0cjLq7p/4ymsl/yzPuBmJXDAPLfi
e+54mcew44Pji0pOjHfFI15zHlxbr8I/d5r58WLepjdA10dlqV3xMQyZSwtrvDgz
PHPGbishGhNcCDKozA6Nhb3Z83XUekL7tTlAjfQTMFnCVfwF41h32C9KyVwnTw9J
Gabknw/01ezvDoMsLHRq0efxHDFuYFt24/sKiE3DB5ikpZwH++wLrK16yd6/zAh9
4FTDgHlKiAmsCKjdXQeL4cFCd6xhSl+oojD/lRTGJ2c6c5dAxYAOTaZ15EvCbpxm
zC0R/WTAhcNFFe9wlPDdYvYOYtrA7JJ3R06hyjojJ5JbOJ9iSUJPrOFQZgt7Zzwi
oyxxgFGJF60tbgpqZEH55HHnvUtchzUoUR+Q0M9R9qp7mDPPio8mCcLcMXLYXRnM
IzibHu1unCgN3rcOfrVZu9IK+oSwNdvpA1slTcwT3jcWlnZRVaJEEfpl2kbf0iFO
vTxOrE+vP5omDrFtbJ4otiGFbd9Rdb0OE6rupLFr7gAuRVv8uBgeXT+rt8xdEt3o
LoY0lGn5qqLRk17r24GzBFT6LnuMUR2AyVPTRm7nOcMHIsf2PAIEVSHDs59FSLIv
UD2Ecgv9FM1xFlVP2/qMfC+ozQXCYytleqSZkuvRB3wxWjo3/6x15x2Gtux7zxEt
1NS9QL9Ie4ctx/fI887ks74AAIr5b3Yf4Ohy1qL21Djtme+Y46HwiM+0NhEXpN++
ao34chc1RxuXukfZxafO2YwVRws+OYRT96/8JAi2RPHqMbMJhFMas6mRrn0CCpUZ
xiS/haN49eR5kxKhr5nkAvbNvNOiiyfUOQWOJm2OFYn3e3xxZ6dA4MysGK4hf1VE
6RF50ssyDFEwWrDCN+b9KTJ7/OmqL4cLxNgrdLICLjexqtc2Y2Hjy/nCRBXiP0qL
Xacmp5b3myRkLhPMKsDGgWl9QNRbDKXeLQAeq8nb6D8dtEdjour0l8r8JfPvM5Yy
PisIGXlhrWZC44edJJYkui7DIIGWEyL4Vi/QUCebfeXFQQC/DepDai1fNNuLh4kI
b/dbcZuQttRtevPRxQfsZicgtz5CQQ69fa1SRW0smLY5rRTkAI2q7vP2oUdDAObQ
uFUn3zri1Ri0hFFnvNPLrd4fR8r3W9pDyQy2u3LG0jMUmNYRAL8ui1cpx6IAuEWF
HCo3tNULgFWgzm7pWC9pNPhw1kr/HIqUX/49gu8o+11kZ6dA9irdz5ioxPDAPEFj
nC1fR8SElKAR55Qq3o04MMYWqHWXpphhKBsZKclkoJmrngClo9gavWli/oDk719X
Tat3c1pI4S5f7hwxsy2Hfpqh93+vgIlJUwHvygYyh4BAWOWqlTuy6CCRFW7nB/Wr
6jpZUGECR1EdH6cCEFcoeSkvDFyJBzHvRQ95V4PtVKJeQuKVkwu6xJuVITwqtIeB
nrJzah2K+NAQFqa1mEnl236yfXYKP0e3j5ioBpr+kK2Gb6P4x2DjwPxqK3qv90wy
AwsXopaxgjJ1K6N5YagEwxTwq2iPXljRWpzBXFv5p8x0r8cyIJXJuIywcqZjegn4
ryIGxCpQDU+juMvM83UW+24F6Bau0vWaY0PdSVrx3/gnuXwjZCB0l6H+K/CrAieH
8fxtAGOpjydBUiEnKLiSsYL/rzfIg8bhQtt6p7IEEhznsFABpYZ6I0PU9YEbPJbW
+SkWkUAn5TlPZ0UURrwnfO6264O7VegzkJKT2FnXrueEWFkF9w7UrNM49KqpZaIK
onYRdoH9bUHZj7yIyMYcntWCUm92/ft8oHrM6hIpwGeoq2kR2cTQZPG+vOkDpc4C
XF6ULhRoohncbV1Nq9kQ5WfVmB575aBpb+t0ezf773AjXw1ZcJgsvMpexCuKZ0aN
YeaZjpy0IRzmS3kAG08PmeWaSmNZ5UsgpcE98UD82Rw3h4OK+P0njFcvuS5kXiJ9
fYk/KIrDX0gQ1zLV7MZGzn1Q1SWjSx7ZZ4EnQufYGyr9oCULYBcg7271kVHihgcI
jhClKUm2ntDd4d0ULeu8f4UKp3w0yW1Z8g8ZtGFaSE4WgnM8xXZBIHvh4Lwpekjt
MfTCH04w3lpd8WfyYUfIHxSQSRJQdQIXGJrWluNrpkd6aKK5ZfXPa37NhTIV786s
BTJqFqjYqDCviaIXP0JFCEetnpXnq5NAUv8nUr5aMyNmSmOhQY+cWH2FXZdJKIMv
uCSizOyPQHIc5GUoIxGkkpXNepeODGBw1C9lglB3TpBkcD3JVl//JomWEgzbtVg7
FrWusPyWipkPlJ0vDwD8bXNdfjBEkwEQb8y1doqY5ig0dnSxsN5PcB4W6Q7ODvvc
b8ivGeJr3IwwxvekV3L9/nITgiw3pIU+WAcZHQMfAmrekuL1iRhwP54pGY7m2ZBC
57Tn1tUELubZ/pTRkYjaFJ2MwiCNWDcor4SiCqlqM8tR0sOmqg9Vcx191Bu0n7su
9izcDv00Kgywtj4WhUe6iaAJBT+D/AiEKcERYp3bQdiHZpFrShOyaBxjhw7MoHIV
zLyvDDvnE8a0BKW6dvGRmwcnrva17ZwwI4XJxKtpRiL8+/TtTFF5NEn3ZiMMBKyf
efeQ60oglDtrUNdWdRCeICdI7EJIiEto1dm0sFgkZC3Ykr1wpokDxs4wqDci7OjH
ne3ECUeG/994ABZVbJPdf/cQEKpNhXiDoYKQf/7Ms0fhrrHiFkVOvvXIlY3y4Vbh
vGItP3L9PKouVIQDrUOk+tPAjUtpCGL88RLlBNM1Q0xOTZdu4gLBUMLoXgkEur+7
ssRRbXjB2RKq8VDMy+io9zR/GWFtXYoBPKvVd4ZgAisfx8LFIiOFSmG/IiCyLemb
0k6h27xXepDBz/xhe0r7JQCyMuP7cKwASiNrM/zrck5aOhynJ1Fiyep1VE5pY6LO
1vQUy7adtttYEibhBYZU0AQzG1/agwRoDWdkEhiLrUMdMv8GpWeP8dlFSre0CPu1
q2bgh2wVOhOZ8oew7ABBJU9elgZC1pVz4d6gHxCiADAge4rDqc4D23hCHVSp5mgo
RT7wgWnlRCkiuMcm/pGH/SZ11jOYxp5BkLZONyJzGz8Wgp76H7FH10/CCdI+BuVW
7Dd3vyqd9FZwRzmxbOZ0gx2iyeahhTMbS3ttfN3cF5pUNpW626SgIJ2LC482MNAv
iPcxYs371scp6O6GaJlgt9R9lnwTGI24nI1v2M2gySf9Rofxvj0lIKxR1URN3Zd0
ke3g0NciufhCCwNxDeTvOw4C/kQB7kYi/FHjXo2chSW/djhCW9kcoKVW6PNoI0VK
1DPDHZjHwNDTktQPI7NvwKFg57BpGJoP7jcjv24BvHjO1nKwgkzSLPj+u+H1/Zg1
jaee96gZUKSBvAFGUeOAq045/BCGtvAwRKKgnBGtpuZM+wBNCW7yfeDGsUANEdB3
tv/LJPBArHTmNF4yoreHDGj3UyDA+9dy34S0PoEVlnUAc1YEp8KzYZDOlicX72i2
6Gdiak4wRRq2L6wLD6HS4mEfNJh8AjiwCLEronP6NlK3mGBjWJjYPnCRzzzhu/PI
jjNQkDn0b+W52Od3vAaWZAefDqVjS8+XeWKVLT7GCxPgxj+1cBCPUUwV5zAUNMsX
JarORx/eLwwYJpZuE67xvQurdEnX45l8T3hh9FZo0zlrigmVuDcBOJ09vJtTVf5G
TxB+RWGTidMRKE8kSU8GHyBgw8FBWJxLMwfh5RlTuD8Xyvfi1m8chWbD/J/c/Kwy
E3a1I9Ey7ZprTnv7b0UXaw9DE8VlcQVe3I+2OjwjRzlRBun8AuFESb5kNNI4p53d
6zer2SeVuqihv0L7TyzMVqdPwkAmJKmlC8U9cHXJPpxdD2RBe/cojQLjX5hTckoF
MY3s3E+S18DB7CjfJ5k54QgRkRDnsJvkD+Im32jz8izk+i6mhwAnmdkbb3oh1Ttu
v+Za3yr+fIhImdpPMeyN2/R9n++6Y22MblaR3+vBXgdbvmPwp5Lr09BxxJWHiwv7
EBQHZEtBNUXWstoGkT/6W0MU8IJxM3s9ih8uxaQBb3mXRtWOnmpBCePW+nVv2LV/
sLS6b8wFjNrLXJ65BQfhO+prBGoH930vWXu7WX5KHLC2X7qtd9YM6/IWM50SOV/M
sTdzfwNwDh/9ok3092o8moem8MXxxc5zBJVYfOYcFLfMytqOHZSnbSm10aBsFFiX
vBH9ZLbHR/GLsXftgx+OUDhXeUWGIXPiWXBDgkP8N8uPJiEygNYWKGGoB0MTo38B
5iFDQNh3kcQ6C4nMqjFYyMsgMJPJb/aSSYguMuMmNI9PML7XMtrieqPU0LCn/OU3
UpM12fAm21ic6oQobBmpRjA2eYuXwYf0Sh2P6cqM9VkSiEWit5VCs3d8Nc9F+W26
pzgVSdN8WXCy2B2jBAAkJZBiQpoYZq/ee+A5m8WhnAlqCvHvW3qo9MplNNO3JDQP
n1a88PcBBYI0oadOwOLz118JZM7NgcLvp1Dl4i2Ckvo1ZjPuXF+4UEpTRXVb5nCR
fpOtJj40Btb3AzELA2GiWGITrS/hFUgy7JBitWzrmw0pe7OMepaWxLyq8Va7UTx9
Fm0lmlPPZqW1NBYRIpZyLq+ZO2GaDabYSpbBtJymExIiQFnamtNcsEmDobXYOyEi
lC6+nVgOJywiMuVHdoKU/EPAL8JhZbsfX1bj7rah3YQ0bsAEjoym0IfRUZDCDwr0
+QplYQai+0I8XolQ1Vz0nsChJ16iQEDkdo/1RTQUdqR+cOuZ+xTag02rY0aEqe58
5RMfQUy9j+P/m7wp3Q1LUbA/yO2/4XcjdOW8UtN9RXacEnct2P4w13LSIzIFtTwt
G2w6yWdEiQetyT6/ZRKcvcXWO/Zw6dGsuH962IdOob0cRfrEOu9TANm0B0wGa7e3
G1JqhKIOsYU1RtTx5xRSQ/Hzp9quYCBYFui68Zk6qer4m7o4TedzPUWeUHqmNnle
Id8I/6fnqKb1VdmGRat6WTmmTwpNMgxJ5IttTALEq8LqNQVqMeq/A8s112+6ADPv
4aqSTOdAg3EbLVCRz7Mggmw4gL82V5/o2uYylFhALJlDTioRGPi3iEZygoVLCsvT
IkHcFjw+zZxVZ3qH2sb0JuzFSL/bkCMgD4oAWf67O2fpV8+PjWN5907KITwCw2Qz
qnI6dMDGYNIAaC8VWvtXjUu3D7zK1s0BYIoch9n3F74vuRc+YFIsB4a3dIywyvxw
vbr0KXlmBhSmWr3IMBBk/WI81JLGz9BsORuQT9f1YzKRG5L7lMynsPIb6XlJc4oc
YD2lOxcaMDFsZKxWr/Q55RMelTkmuJmO/RcvClDy3tNWU1asDkPl7QncIt8jEo7w
ZtihJUD25EblwE7kJrLFFW3h2jYN8EixQpS8vvSPYk/OxDkhsqalxTOtG7bBXK8I
DhVpG1cWyFfyziygNZ9zJeexnz3/lHrxbsFienxn9pifb2X8YgJZW/ewy8mER2Bj
fraVn2ULpJrbk7zWXFK405niOg9yAzV0Zaxr7lsv6Z4bsKT056Peq6moYBclZwMy
KzBNxXZ6NL27Vuc7BziVRwhZ7ycqJXv1D9s73A0XzSe+AStPrkl5qT4G7cnghvGu
AfM/XkLfIM0vBEXWwxnSk07fYXxPRT3Fmp9qKT5tHkg2eXtoB7+4oazP7Tdy5YZd
QlInOa6Zg1ues2JpYnnMV1yEv7j3zIpPiP5gkf2YG9NRO9Z7bsMhF4e721+tVDHU
9BOv1B7RktnTzzHAMtEoi+Zh+5teS07XEAgjgPjeerqIFxn7dr0BjhxO5AsplzGu
haBnAQLw6BnwW88rDfAFupd0eEVvaKNTdEo+TovR9SHhhKfseT2umQ6fwC2IB0VG
epI1dImc8rK9p7ipS0c+v/PUhodxOJmXY7LHYab82RmPgOADxzU+A/ESWcwhVlCO
1HY3gG37hO1wY2fGPVL5vvaAOMQGXVxWlWFfSW4zgP7E/QHcQ0A/9F6DwUJoT0zF
4CiqEnRSRF1ABOpkdKKgqfif7Jthp2uxpNos7REpoRC2ztGv+3GTSWUE1O57oZiV
RR2rxTSv5zQ8jXmhVhOlVFAy2BUsWtf/4NKfJcAQsAsEUf1eiBgKbwoG7Mp3HKHR
/FKF1mHAhyf1Vk66Y6ySEyWFwabs32NGmSczMYoESXpJUyUK4YGGMag+Xem5mMLt
zXftIzibQD2o30WJzChWLO+Zkuax6c8NzdcHydEJLkoKps0svwqiXHt/xSnbyh1d
y9awbRBrVl3/zVAlZAxesbTTGLcpGAeWKa5M09TBkanDPOc6SmrSdlMPbdHPokP5
lBEtK9XBDkUNp5KQgn1E9knQxuDtSoOyWnFOBJV3ippyKx/nsdfRxr1Gt2WGzksf
QUGFXvsUVzKZ2fpw9LDKzUBjG80gQrkAxAqgAEs4SlBC1S0q7eVOItXUdzO5Pu6a
V7KvJ+hAmzuln522WHaMXPBCy6hhuhED3XD03KvrT77gouVXNRQmaP1Mzy4sp49/
LVS+yHL6ckHa+0hUfWels5qi7g2YzyZJTNP5zXC6I7YdPYnO8jWHWDcTFFt36CiF
7W3f42VHVxi6u/yIaxntXjMEvErzpzELV1TvnP+dBYioMOGocbUak5/qnjYhThw+
BdGjriSBc6XUZq1Rf/gp18Bz1i0ngY468axyxay8q4f09jEYVbkDptcDdbm5jegW
kTW1Yv2mZb1pgcg7zJaFnZWP+Q7zr2OdzZqHiYd1kpOPDoccS3YxN32DigYv/koM
QewnwSNag/vW4OQivysUi5MK0WzgKldbgTzstkHQ1WLfpFroVxSnxSl0PufQ32g6
xkmphP/iTvyhPALArNc0cjRB0d2SzA+NdnuEavczy07IpN8NUyzThVzg+hUEA4En
Nq0c3Ph3h851zqlygMItJYj7mv1plNYqghW64N54jdNN8UqOjbt5PNqPAMwGcmWQ
FBj35GEoPvdoClzRXNKgGuivt/ZXEzqVeh6QYvtUtjfEik5D0GM97ZdNl7zD3N9n
sUrEC32w33VuXJjOsr7HFR6olHu6xRErcNDn7DyRfZ0pA3zbMdFWfSAcZYqdYUrd
Xafp+u2IAd9Wp3AM2g9X9FPx9APuTPPrK0oO+zBgez/UuWNqkplB2xEbBRM5XC5A
WbWyRtc/U0MWPOn1RiL2Hhgf4yAPFmCXwg9D5ox+OI1aD+nQBHyfAN/nABaNqUt2
iV9Ii0vM8pxltqKJ/mQXnq5W1s/AV3ajDjXRnwzBKQBn9b8GeoNI74RkCQiF6vyR
DQgDzYNSgDWI2G6k78MNvdlbXyAGzyHDZolbMAQvT4sZp6i9RJmk0w40T+uMohSf
PC/TsbWD6QuNeFYBIupWNiOj57zwOzA4IS23rZc6M4eokXzC82LJZj92aNfqm5Od
QCMEpPCKoMfi84hhe6AQE5+aOyvaL37eeuXEU3h0xnFp95myXMa13L7HeqMyCNTj
9njKDtvfV7WjRNdZGlApioN4s++2hXTgZauZQ9ir6X7eOKHynnFvA+2z6FOFR85a
N/dDlBuJGYZn1kIMjpHfTDPUYXoAf3CBwbwK2+nRmVAvePKCW++hVIoFt8kb8wDT
2CDc781/MvnDOHF94sJnpjpcjlcugnS0taaQYhItbsMxfyE8gi4viAhcwMzp5c2R
YoBHi8zyZ1scQZgUA/wCHdkNMci92laAk2AEoGPXmGZYKHytRbeQWYvkmcH70VMH
chxYFdA18sIEKPk+sB1TwMLbU+GzGDY1p/LAY0RZyR4aYJKVc8MurzsF5E5d+pqx
tehEqESt1WM4gQtd6w4Qqarf8pFuFqy1GxBooC4vzUIMCkfxMjbTNEA01VBzFHSp
roYDzJLRGHqgbN5ctC6eJ57sMt3JtsbDHWK3TgybOSxZbjBUSrR7zYgZfo8YoiDx
YlFw8wwNxQgZP5nPzMPpEXwU1SBNahzxEL6zZ3tDmmF9xpWRgU/uz7g0SSYahgXg
aM50VfL7XKgkdEnY1Mu2JtQvj5D0Fys1LSr/9tztSIaFa2UBjO0nZgYhs2lloD3H
0PuXeT6hu+ypcr1fIFQZVTH0W1vBxLpqNTIe4I0Hq0AA1f8R9SGb1DrM9BmjCy90
rBAEx0RESsiQw7cKVTqjoGAWMLXTUshtriFIc9+Q6SjYWcMcSC8uLZQrihdphByi
13kNVN7OvVDSj44OD/DCltKyE9zI+D4xbaZAE9HbDpTxqQzy/A86pHzLQspj16yN
t7q8nv4tlRdPZOFb2snpoJVn9IG9ncRbPHPvOhibXvAnGHeeRzyBdZ6eOx7PfjU2
3/Kxwb4NuoXT827Zc89/1oCnJ1QfitLMzwKuOlPKXtdAsi++dpmrNuADNXhdrF1/
gNjN9r8FQTo2YqPqDD0w+wPIR6IzDEh6/+Pq6rlh/JPGiC3b2CRcm08idm2HkU/R
GWBLgDaePyoAwdZzkSWQT5KFYl0FVpc9uVa+DeTuHwUMgj9KXMvaQWI7LILBR/qH
itP+AjBjpTIyalKsknvkUVj0rjhBg5VGLHqP4t6oHnylDeE+//llPYwGbWdl0+sy
dfE+npaoGc87se6ZaVmW/yFvZms9S5jBr73j8IL1KTK7pmof+VkmSw5DNdM52NaP
k0RVJY/DDrVKr+ubNkVv+suYnNK/CqfF0Bx0G4LqfyJjakAijoLKTVBpIKCdV0s4
RTm7x5GBH+hZGBHS7ZEiMQ3VAdGo1j6aWCsG1i9Y7HnqEfvqhYKNn5iuNRuu+XQm
AGuzfgIsGQWt/xAjz+4H6q3SyMXPHdqyE5UCzY+mmnVB15O8O9m592Iv2e3iAAP1
Y/TApd5+hdry/N32B5cHNisrxNqR2QkjApgdNGIUZLKXsD0eHO3GdVLNL2Hn8Tq/
p2kSGe4BpjrOE2t345R5acMWh00BOtrJBBu26Bniw0PgOaAMm5UqdUAhKM/CXbkX
bKwnoSJlhe57eZO1C33EJpYJRyaGpH7K3Dhsd4fIyh31Jlpa1MAxxSXvZorqqJtn
EIUcgFdoxSth6kZGag7yY/Zi/95aeDkRJo6fNmlofAq7cDDsTAPU+vetCqXmZJn2
Fo7OiwHNcKE37ZI46DTobg==
`pragma protect end_protected
