`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="galaxsim"
`pragma protect encrypt_agent_info="https://www.x-epic.com"
`pragma protect key_keyowner="x-epic"
`pragma protect key_keyname="rsa-key1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
w/uBVGAqA9GnKHlxeVRad8/df9Ty4f9jtGD/GseiJCH1SLfEY8dIXIKZH8ez4wmW
sgEuOuYLsCE8S4dMRlCch/Dl/pondbfn/CuR9BUM5gmg9mPPVj2iyJV2lB/gK9/N
+BB1QxV3oJcEZD5v5ywfiY34y47xZUp1VI+1s345i8SG8MjljR5wx7iwoclni8GZ
WgublJBugHpVJHqw+kFUcxO1siWIwHTOHNbYXYYdL0WWVQGSGq6bs7dTSatz1dpG
b46I/uBbylH9Mp64m4opsVdcO/G0Tw9LT1K+4ShCfz1QyMfr8zdvolAm1n4m5wBx
66tv5bB+00Wc1SdY+0EybQ==
`pragma protect key_keyowner="Xilinx"
`pragma protect key_keyname="xilinxt_2019_02"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
h61tEHkC52n0CbUulugQC6rUKjaZ91QV3N6nmZT3hze4QutyUkvIsvQsABssVo4J
VrlAW0I1vqLc9gd0Y1cgFzsmzEGYqe8c7v7ew4nQ7Md8pNC1c9M0x6XsM65HPXzx
/w5+ckYCvPMZdZfctVi0fglvQqYW+pYPAySkeB6ZUhlD0dnJb6thr02UGySQkGn0
Cdv04v2InqLfwUrO5PpnM/K8PpOoQppFZS2KRyMOACmzgpkqztuGdwzukudjLafb
ZXpifHQNCwmHDnOkCQM5iyzwA2o0krDSIYoNmLt8kGD+a4Dp7w/yiAsyavMhpOfh
1UkPZAENXyejg+n79pX+dA==
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`pragma protect key_block
r+nEl55QG2zbJ44mRECeGRrcxuEu8glDTezQM+lrEMv6BcEPeaguMetTIsBSX+ls
lZtPrTvcxKuVaeUNN35xTsgKaOf8m4DF1m0VzORQCHjRACp1b7aeodei+yfzH7sr
rLmvROKxfttbc4mQKkoz7teFlsFZnMarlytvFPqNfgE=
`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
hLLPLlDoTl0iyCi2YLu8ZSi7HG+wEuf0rX9j6V4mwcKiNAr/iEHGSvuU9R3zcNKc
bdRApFtbuUyibIecjVl4UCjXPUzEwNjVSKzDPhMeME3W9gNZUjxRtOB1HR0dDHDc
oxVK4CiX0qaBc7VvwiGTYQL6/od8bDSGfvCwyVG7sFGC9rc8+tZNDRvItnmYtm5w
I/RbRXCspQbbtkxBXouNv5o3nFgPQboIl6VhpQVKDo8KSHalqSXXB3454wepKHyE
p9O1g2l/bWZ0ev60fnKsuZ89rY2JapkuUb4eawhXCWqCjMk3J0AngOozHinHS1Jd
wX6WFwvXVLwDFYgTLE4Q0w==
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP15_1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
H5wtnhhNUqyg0RYwSH2Znx7Dns/JxNak1HyLvX5M992+aYYw8pFuVPtNh2QGpZfe
H4iWSR8NCR4r+1SZibWLQr+UfT0kqW7Lo9Tqi/4bbGhKHRSfrf/WqpeJqOm2E/cb
zdYCbW3s6pzA4fT1SbW8VLo20avI8uP+nH1kBhxommFBmbRx1L7q9QZV13sfiTVn
dSlzUasGjm2vcQMIMh5b5DcYfj4usLBzVslA1To14jxlyRrmqzUBOAdLJg3hF3/i
maK1JD4FCQICEeuRdJX/91KUg+l3nnxEMaiWNLMP+X8e6seMEXiwndPv9gBGTplJ
xW2U1xwO4gtqYU2wHPuw3g==

`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 7952)
`pragma protect data_block
IfyNkEPPEdoBMK9oenYtPec2ftmLVzKBUUoqCF5oIvjFsniBy9Yvhu7qsmfx+k5c
j+1XQCoTC3B3jxp2+HR4GRu2i8MTq+rKPTXRahQNOU1C9441eaSPAHcchgaRP272
EfM5GprzPyRpixsuEv990K9qyrVav/1FyM3wvCUBfKA0HSb5RhH1dtG/xIkbk7jm
opvBBNhyPpfxKaQ+fy2A20bY033BHi1HJC+VG6e/n+2sSwWGVkMDzXsvLHhTwDZZ
mnGyLuoTgYpsA19qdi4cqi/Cp/fk9RLjy/eWwktmFYNFGq7CmfZKwlotD9Emhmrk
YRqNbIO8hi0wf9J4nL984geu/5XklqfqpRZanUol2fcUwJhJbvgIV7Oelq3gnlVB
mbsacLz34ibqUzjGFJVUW/Q6wyOm+SDGdIgaGVudodv4N+m1e1nrA6EXkC7HApj4
6xOx2LAQRTnXBWuB57DWxRIb1SZvFBXd9IlGCckFX/9mnmtv1I3XnCZEa7vkQuo8
3ScSLM4w6kG38r5KVMMw0poZlFDSRsYAFxW7tK0gFkgQOdmVsXv5SeyitYMDYrhi
2D66hXyuPQx9LkdRfrkkarU18bds6yF/ifukV5+z25vJd42oh7xPT+dwTLo4kJtX
FPzcwzvMZnbB8OhUYYF9ZkQKc1nZ1lCiTxz/9lHeNnfFRL+1xFCKe4g2UZ6LW1ko
iDvc9n5VP1oS6OMR26wdWc8CuHv7rbYnTRr/9MmTdsHVNEhJzoEWqXO3fet6xw4H
S3sn7KwwQLrbG7m3/42tBNGfYXO9Wns2C+Nn3rleYt6H89lTyPeoB7S5M+mfMuWB
vigc9H/2bdQcE6tX7ysMQd9g/vz8UXSK8syTa165dNwbdXeBefNDtkgVdfpGmMtP
B1R7qJyONQK2AsoKDQpgOXf13i2FQxdDBvnWiDwQLKkE2YukEsbQMm/mOhBZ7K1+
5V1jI2uJitQUCnCvdRFAlC0YM4sCAIF3F8N1gk2AkpEPj6QZOEXSNIqC4VtERkpm
w1chJnPsK7SVoTxAaSrE8zBUvO4Pq82VbHzyMEyi9pRUpxt0c4kguPnsFRtnDojO
cM210yE0bRjxZM1keXEzRhtYoiw/BjZkOUkhrW49M1lOety9MmGEnRtWnB64tEIp
i47gppQOkZtoNd6Iu0ZrmQl0Xnr1MHhyFV63ZDA/dKyoD6frmLgTse7SVucP+pnO
8E7Z9qN7E289EGxVNlPG2+cJtD03jh2Q+kzcbvVdORA3pit1oH3NabWkREpJT0a/
EBtuzZUbJv8wKEq+AqEPu5jBMKc7S09xNgt/4dxPzI6mIOOzLWihrf7QlQKJAOOB
qz40nqDcYM6Ljh0WCQcYPxAIp0lk2IbaQD3gw9n3HsJy753SpJBQ1OTe6z7xgwVt
DzM845fJRZUxkcYrcoekpaUvjrSVURfIyLGkZ0Hzq4vzVR7OLpFQJn/mPN7U2Pz5
WegTLW+6c1ymGGKLGMNl8OH+N3JwWQC5bFAtHczOoFXf4kWOfxm0Hv8yadc43TzZ
l2XwuL+DSY1t0X1HBcNrDW2WcBsScIOmZ6/jGor7+NQztEVeH5mB98un1mAnbfmd
ooAAoAmioIE5v4YC+lfJm82548HkA10oKjOdvYShJrSqSBqPZzXN/bgKI6VzleSg
XperFg1hWSJx1Q4XipGUY7Wjtra7/iFxUBkVzFGTFuhFX5t674tJkfqcF33evKce
ES5uCBD351V8agXMlKNQxy13Oc8cf4dmoUKsU34HyLwwVQJaQmwZCy+xVpF5EYyy
IyvrRt3EYhu+CvbsxNZncbOygUrh+sAp5NyixZvm/sZWi+AnUom6TLTjZCmwr6g0
UwBvihfCqsTTJrbIiNcJnbtZOBLKqgPKO4NGC4d3HOLOVZykR9MJTpYbR5NMRuTt
MfpQXTidaFc+ZkqWXv/cspO4eI3S8EMQSBF4Mv8rSEv5SQo1l4En2tJDB1dOsSqr
vej3W+lX1zFeur+bqBsCM35hU6eiq8IpUhlLueQdmXbUTze9ZrmKccAzyAbqOHNc
TswrDu0F2oFerGGZz4fRjSFLgKwN7P+9cp1AkEbBak1Fe7Lfsse77J3VI3npAv6k
1YMGLY1OtmpZTdAJnb/2dLK0XHoFozUxeAvRXJIBWSvJCn/AqvoiCut+syy1JR2q
7aTYXxroSA1iIj9DisvOQ2JsjYyLZIAYSc7/NfFIZ8ufsr+8VCDF9eirkCsfuHSy
yVDjFcqY+tEZqd2OcXs5ZKr0Wo1RoFG0zQ4jZ0c67fLf5Ho2WQiGkvsdCrtOU6FX
m4dUj7Hf3s0sbI5Xntb0Dk0cY2LpDdGg1quC0N64Lx7Wjfi7UKPUQJhkooHzZ9AW
6RTHDwZyQxp9x+jnDaMpElCqJczJK0ndvL2DrH8guV6ctNrYGxjxoPKltdzqdTam
TxoAK6tTEsEAsB+2J3815DyGf8oKT//9uAn3T27rQckvxvfW0fZeB7m54gF804Fe
WWTpa2kme5aMsZ/gwMP4jkPmPiypj0x6Ae+XWYqqd8WL0sqnOrqn3ESWiKylZGqg
v7IHfpWQAhiVgaMnY8xMhL0qHZcRt2/hbtizFzbZCXy8ryZcr+BS8uho4QU+NXFR
stzU7EoNWZuvbun/pOy6B67oU5D2gxKEPKAKtTKDP2y8//4QOVb5FCWRWS/NecKM
2xcD5MwvMQpMFzU1eBVjkduL8E7VgfYn9e6vBwabXSiDFrRbaEJ0AvRe/Hk1vm/E
49Xj0MQ/FF43i0X6DXFWA3wPiTQdPOP3rTRor4FyvT878EFrNBscps3pgx3aWNZO
4HTLEaLlt23PQwBtb+BS8019vTIeTsst9sH/VAZXmCQg0R2pTK+ByerLcVt6Xnxs
HGEzX6WZsXk1lnzL7i0GCsLcqEioeowcgk82pbFZjrysJMpfpoQ5ScFY6+gktaT2
DIoYEj7KWWQ2RIiGnL3upmZlypy6EVL21HEGGfB5YlTOulIYd4+PkGJaI+P9pIqH
pgmckEr4F32hiYyOdrrZxeDyXALCITqWJv32wc9TJn19t874clJcSnvV/0QfDevK
OdT/yGAwqJaJKsiSJlV1Q2ey+LdwaOtlkWaENu0zjUTOwoeRT3K6shYuZ9e0wNB7
3HjiTMQoJKqPBnhqw9Edm+hybXhq2aj67E/09WpyUlw1IS8OpRsC7TrF0Bln/Shv
xqSJ31mpcp5guun12KSrKAyUaEKK8FP5NLEcMvWEjAA1ECmIYKOuY1ddZSrWJFCG
ZKGsLjZjdro0HNKJO3M+b4Oy9QJy52KU2zOupX1sAQQGkRjCcqtAAFhpouJAZPOa
SxJcrq39+VwPxliIyRnHD5tffgEOpyRfjALD67cZhTzyshu0UOH+zwn8nFRb9d1c
rLAeVudBi/gBEgKt95aSqleKwW5nLARKRi8CNIB2Is0DD3D2zrZSxZ/jT9lIR3o8
GiNr0PbJzi5rnusNYP9ABCUyZ/QJQcQCi3l53U5OttA3uGsExcGlqOsUBb92TMLg
TLPkL4ai/8U/wJ1EyFq9GG790DvPM2XmI0RdzNks36MJeONGNUeCGzl9vuNYKQ3e
LiN4KzUAmTX/e0BocuGO8LmLQPktNHLbYlPgtKHTb19PlCOF2/qxFOKgutg6FiWm
PRqaPbehIgo91yqqoGLkA6FAiKmRqqM/3I9xfr5Y4HLrPFNbuWSYEAHirXKfMEh6
stitzWhnoTXEd3UnR5i/ndx12oche7bC3qpV4ihc2uGNpE3D7/RyjX40KOVHESr/
dEZGLJ9uLzbYiWVt+UR2thKIwvlAOMVKVVyb802jWQjqwD4v5eIcTookilFc224K
YUhb9FLWJFXyT2xvrneHUXm7KGVpnfRL+jGVG/n9ynlzo8o93Z4hKrhfh7W61Jwa
ot5vxSxEoicev4XVh/6i3muSAQAvh5yOQY9B6Q2w0l893fPXTgigSKoGlAZFMa16
nSKPDvZMHdltVXMQ3HxG1sw9BoMalXJ507Ffdpr2ueqKjuVOalgwvEh410VPD/1Z
TvPmIH04EL1+e6qRKo+k6L9nptKMpyxM63U/ZUqw7VGs3TmJ6LXTS5Ftx9h+O4S8
JFFydNNJyQ27zU8FvMBjbij+89kMZFJfBFp2zeEGbCB6sK+X5j0TUbiLFXMRIIeM
y08wmX5y99Ez5AJfjzVFNsxI07vE4iEJV+lJ2AIX04RLQFQ4yEDA/aE/c93jNPqW
ncxSD357vIPdAkuXHlHairegQjGvvwnallsK6E8WTrVjKP5/cpcioUHCIVZu4IV/
niO9Qatewpb9iivQ5zLqZmb6HuCre1A6HYGkTayDpcPlNOYCkXei+Kwp3fHIsnTj
JmMNAeUUTa00f4kGOA3bNv6rhsqkUeu4gbcvKZa7SNzJ6WF9gqQEJEx/GpUEjN2Z
7RDXCRbV+mX6EnYyz7iKutDLxtJw0AddnrY8r955vxAfVb9VRwBKwenqXgPc1w46
jYGVzrw+Vd7Dm/fqnNmM611If0jsbGSyLSwjh8NlBfA/8HVswpByHJmpSlsfj048
BJwja5EG14DJxZlVQz1LyL51OGhbWBwY16szWvWEjsVq7+d5hKxHUnnit9LCJ6tx
5N9Vd5FptywiXhK8Ze+7xdMqlbyHfdlslFqzKIgSDq6T6ioBOEFXDMrnoXsfjDsq
siGoOUF5MxD0YPTv0v4gND33auuok3DELaM9m81zRspZs1W098fAs01EsjzNY7RY
xHBEa/3u9XyzA70MF2qKl32fjKlaN6DqQpsgFX7QpNbHfYTfY35An1VLy6abknWb
L1KtQa/ZjsJYiEa5UEn1RVOLXxxsvZ16Bi1c0tMi5YNZIbrsUHvvFVm4DOKmI0qP
dmb925uIp9zDs9oHMxZRaPkt2K6L7jfAJKUEi8GyFTTZD3kYFaFdgPOecoUgSnAq
tVlAH8XHV91YhI1P7mRrNrc9TNPlBiBNN0U47Q3hcvaefjyh2hjdLLGwPnY4+PiZ
0m2k0cpMyC/19bu8/+8c7zHUbjTENKZoTDcE1QysPJTdO7ByY/7ohleP9gDaRcND
j6LLSQN/CJuPe4+P1N5upq4S9WinpRkRRydTffEkspLV6Um/9exO63qwhTigGlMv
1ISInT2oiXj5iWbWv0IK6eyLIIngP3vGI2QulcRgbciz4zeO6DzwowLuC6dOCrOy
IevP+lhPnUZ4kuu4o9KtWjmw8me1IG+A0D9q03TuVcTcn8jQqKYo9f9yi/Hl+Lak
59Rk9iZNxHO/4+IuIWGFM20ys8d0KwY9iys8u23vELKpyTjd+W0Q93jItGgbAo4k
VJNEln00IANc9jQpbOeFszVzcEUX3i+ZKrc5dP4otMsMyAUI1U1x1feGvyKwLGao
HPSDo8wPm46w4CcRPwPAkZcdaFNtEmg6kH/zhuUV9fCqK1OYmU9Ve4ffmKs7WSAH
Pctddmfxgj5QQzZknWkELhBoBUYb5WqR2QRnv2qBANXR9OOwJbaDkNpS2t8E9QN/
g8zmv+aIAJrtr109OEiXqlD1wFaVgTO3lOEz7xUbhQZURE3m9gdPb0CBqT1ACA95
1t7+MPtykJaG5L6bVSTaYPYZAsNCI6ZX95ORwTdlvTA4qKaBp1tg0sNtinQTBsn5
2vQ3S9sQvoTTr92Xe+vZYRQrVTDgKh2uRK60rT9KsbIBPWCnAI0K/72FssyKrb8M
d9daoxd9AMlBBnpOYfcTg5jWe/5dkU+1CNAw2HRojwaLW5YM6vYLi5Nmzi51z+ZW
jhZS5AsML31BWCMMF2JA9vV2Uez2h3GtPem2dcU82hWH2S3WegL2hTVBYmW5frHY
G3qNXiT8lIGm0Fsi2TCesd1XijMH59FR8oUfFIrmyaLkCbsY5LrU1OQz0X2ThihD
9H+u3l4s8DvgXZy0yelX6uI4CwfzE4P0xWIgfVI65lS8vJfZLyAVH3pRGG36Y/se
bn6WeX1Yii/umhdKk0W6Pq+bOUXoZ1gKCM1A1ZqLP61f0DMzKRRBHI005NphU61v
Olf6wB/u6y6wk8t/mQd8o4eximYLxdial6f0stzrPPVJMhqHdhZ9hlE5dHVlre7U
Ot160mlDxlpcT4NpxL1LlXbBAlNUv+7Dqkly9z6di0tszv37kPUOUtUTxwMlhiEX
i5fPO+PSDWRYcX0xtkkP8Y/uEg5WU8LOwRkbVhu/5GWEZK567nMVoq4euwbJVqfw
mcgCiaICaepgjwz5/u0/7w57S0v5cfJy9zTDlmQmOvsf998r5RV/2ab3apUIIryQ
/NdC/krrVm6Amq+MUl1aD6EJqg5iUswNmT2dapTg4BJ/ASkRJW8PdlgyOoA9wUYH
kLizszZIpfVApjat8/ma2aMY5Kl69uy20OlyKtg+Aw6QVSvWUMl7/hRHo3DP4FSI
7u5sCb2hunDSb4lc1au/8WdyfCs1Q6DCAG5/5T0hr3EGXDFIgoVmQLmnFWyaH7Me
pYPDTADdu6dO98QukiaMed3+JXbWQ7IidDHMNpS4wh2qtD+PBJG2AuQriMcW+E2B
Zsue+TdftNo3RFVVFv8RILvjz+LNMhQAnwoVScgekBcImS+iJOYfSSvNc0oRVrGb
eoZcQtYlc61kn7iEiMttbIt/movjmkiWL63efIwetRVLIsF7jKmg6LXWYuhn5dWH
nDzqi2m3L6PmeMmqR3cyj0Hd8QeqoF1FF1B3EBHfKgPsGVout7fupef3ZqXwh0mv
0ZL9bzNMnG6A+qxfMLngpnxywJT7o9jyiR30yoYgBAFbpcG1JNoM56wI265X169e
GxAzMK00/RmiY7ZrSb6ng6vbqXQVu/+51L6Tny1dzDlkgDollnMosrxdrC8Veuxk
5jy4ottF5lMkeF8jyD8ImWRRgrXU0pKiQE1S0c+98h21UST6AO7q0/50GaKrawYe
95hiFwSrAKdWF8Uz0D7goB9lbj735V1MmSlIR/3xrasc2UIcPj3ZHPDdUxxXFeHh
lzRziNpw3s0JdCHjRdSH7akERO47b5ZsPTNKJjvmX4Khlqr5XjQXymkB505GqR69
+aontLUKLUqakljksu8VZ1d83hw22/KjIjoBoH5b+m6TU07tjZUAOZSrQY6cp96y
VLC5ti2UrKKCLhEZngooL2d4aOWRrqum6MEinFGda1+JsGFuqgCjPzDMGzhpppMR
9Rrh0eUb3nfmhCnEvsRncYQU40DV1Et/XWGSKIvxEcGs6vQRcjnyX0G7qg60EROm
zTCZbN3RmG6rwpHccx84m6T4cIUJgn/AuBt0WoA+4a9ZlV0pprSc2VGZIo83FrGX
TLJ9UBS5ylG4cdV8Bqex5rV+w2mnQtc865BB1Sqplb8xXqUnnD/bQWdQDy8pK2iV
LLj3FTcoqIk1PQi/+9yumVH6nU9LiUckiosuPLJwj85DqaZRNP7lzGT9n+3TfqRv
pZic4NrdgTXfiM5rgUcKKIn8+p/mFcuVIcTGq+3r3wTPqKY/umiv/QlPHr+B0wu4
pmjQA/WnYNl1bGJZsUYRT05NunQF8z/TLQRcSQjCdwNd7osRSS54UPVxvfWBCmlc
SQQgea07fRXqROD14GvXhgaFcZJFB0QN2/jSGpX1g2lYHubppHa36CzTSiFDkgmc
4v0HWOktrKcL+hTtAt8olhJYS0xvn8iGo0UaJXgqe1HqcxUtF3osqpn/+IONpXQ1
5L5sXJxvlwkUpsaHHptazy6taACRUnvbWxuxw+hhjiWgOZ6Uht3NjnzTOyawc+/r
VOtQlQeFNIkz74SvUVCWaCmP2IhDsYndb9yHg+DGHdc6LY13CryoAIDv0J637eRB
xD9P6arsjlcH3Yw4YOWCnjfyEjJKXtM/wMfvqYUS8RLM6xXLmj8AqBxzyuaB7XKD
WOPHnn5fM2z2qBmJlTUYjYC//aOysXAWfi8E75wrElRabxsLAwSLH8fMDEXOstfx
HxC/UR4aLE0aG+WupHN9p6wV/GSwLsmIUbPZh0imomuM/5cWbGNch+UuhkCcEowT
KXMu/zG8wnvxtT+xXjdghLI5LqeTOyMUZIp9Cr6wXN9HQ4a8e0i8N/2CNK/6AMs2
VlsFkitWDikU4+WHUExGVUjtaQ7rw9oBjyFYUcu89wDMFRp7Wa84zooDXT1HM/FA
VNxMJKZW0pbldsR3OH9GJen9195e+p2CRiEVtz/19b3fR7mxRP1tLi26EHCEALDU
ezwxV5HqjiGEzr7CbX+VmMdrXLv6F8jusg+7fN4AOtn+rRpTPTPzCie9IJ+awomE
BDYo+FgH22DiQv63+I95puaV9M5q1vyz651EvBGuGHJCCtnd48oL7cdgT8SolBte
2pQZYwLy7TwOaW4DNy1y6mKGkPXb0cU51sAD6Gggt6OeAcBN/HjxqmZoRJhSrQs3
t1JTHHqguo0nA1LSLWUyQGQ00J0ApRJ5yFMSf3L8hEAjhr5X0pFNnl2nijUIZywV
uDIyiDIp0regzRbq7hRnQHppiqFE8VfL12T6dHBbvtRXcKUecTidh31g160ZE+F9
YAbbCvo4YnalIIFKygLZifIF++79XFNTYdRKfPm1nixgPCCqYRBtx6rupGCiQ9Zs
Pxw8yZMOr38p/OMdGfoNAY5TxHpGSyWns/ppe0qNW7mDr9QnLG5Fqjt0qBm7Uku+
0cwECdS2Yx21uUbSYEF+8hGl4oa1o/EFC29itEsesyfJTMaod3XCI2G1GCDou7Xd
F7qwoPZCT1dBTHPr4cRSK8a9xUWtX2inpL0ISMSXQ2+fPJzXUSoiO9ljYtyILRAm
e32OZOXpBtJZTEitzM/xCEx13FeGWYICK5MxXCwNs3wuUNdKpZu+42gLwZayUuaQ
7ta1hdSUhlrdpO+u+frteIHi3PbjMSsmYzHWa8zKcWd/WICmlmbQB7zxWqru8Uq8
+vxBQwMGSSc3JQWxGowZGUWhv6tL+OxOXx2sTtodCB9OD41qt3GPoTZ73XDbBfeq
hkMIXv0oHTAmZ42E2v03pZGFYXTBFMx+GhI1Rs/VsUtLI/pMFw9D1R56szyqmQjM
+EUSkAaGWQy/o5unn9NWbKHcleJhJ7g+4I8opQs9R9I4T05qXgrVLlURU3QHvzS4
tEGX2eS5e2sRdo/L9wcEmlO51QRp2L262kkc97U1j8KEbr/nZjY3+o48lIeNOhPf
0naRJZAbH38Ub1ef6byIPoPoD+/4fGKkhZFzxrWR4FUZW/rWKiDPJvjVEnJnaKQ+
jJ+y38bb8EUDVvbvRRMkANuwivSLkvAg77XlKEjaPOpOE2rauRYTOYQmO5h1lUNx
28p9Ei7rlwyq7AoAqiZwKb4LJxOlGaquA8JCI7OIVTfiLjrDcLJ9JCfEmwQRS6D1
8DAC+79Li4TBiyZ/kcbf4rBTZsTvPwYpsswy+LMsbOxM1Qa+k4XrNC1vwDTFh6Oz
P4uVKjd7bV26u+MSSmD1/Kjbl0M2duK6jfvUH80MCx0ZOhhbecPkIMubv+aDzZvD
DCMIB9lKXtnAkdRYLG5YAfVuV6MYFG9lb6/2oFYMNd5ureYHh1sMPhwHMZaQKtaP
1Itkj8ygR0Uh3OCDgKLEGwdNbbIkWNDFn+jKJipbnHX0lIrXCjEZYHeSe5F+zz6r
xFsMlSPnE+bFeATjSFP1Tx8VhouazxNWLvIgLEBtSZAsGVWVRftA86yxAEgoGnzv
ccSimVVJnqpYyGpqfNguSoa93vgmDmkoFhaSWM8kXixOGB033swIE6bkMMYT2hde
xaM3nfsRPSZ5L/XUjC/M+d871bL/3UMlamCn+KgSDdwYS8Ql+l+EbtlVOl0I5hEs
3aU0NWkI0KcjjFH1Rn9opNybiVtxHNDyTdUq1sLgk7vgykIQSCK2Zmbj6dMg/2QZ
xN0Bhnf5xIqQ3h/tA6jvd6uiJiE7Q2woWoWjTqbtXiRUkBPex2f82fyw4NVHaW1q
/k/PwnYgnCriRd/TJ6lPQSIOHS+YpqMiAQDQM2KHrVSoMl9wAJC3iXi4rTB4c6wj
347JAu6MmqY+zP8mz0hajjCoC9ypcA5NQbjpPctcUFhocWXOWabCwUfT7f3OgPBY
epgOtKivDYBR2Wle9sfx4r0cnYT+lxrdaQDZ5rokYKHn/yGYjbpT8z9e+IIydKN/
lv8SLCZrXTE3uVs+0YJo/X6UltXr0T/bI8CR9LCpOvmH4wG2EOAs41pLRTQzh2cz
Yf0GdDzlT5NqLs24guNMJnx1cULMTndx9ASTYI7rPbyHLjiRaUgC6AIVDEav2WfT
TDXdLB8pEJ1tt7sOBRv55IGwnVKViIP8VvlYMFFRFgM9eYhNPbshiOVDWlq9Rz5y
N2lje92UtOrQpNZQIXNiXGDnV/YjuOWf5t2p5Cp9wCoj4p3bYTkCYMIO3pL4W5zx
aZEPRdsnYcJumNlYg7KaagX/X3XITOXhluW+UKSAg/ED7RB0tj+kq8i0Z++lq4ms
HVWo+0xffcAviiGgpW6hnnivGsaUqHQ1zdVHYFwC6onRP4PI0wb9oOyHgYAH9RTZ
2UcSmH3z3qNnAp93l1u7eeFO9vpd1oc3ZiX+hjptLGB8vbq5O3R6JPOFKsdL2C0E
okXS8QEEd+kWF0WDwnuVFcmXKyZ47LmKYB31nn2LHr8=
`pragma protect end_protected
