`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="galaxsim"
`pragma protect encrypt_agent_info="https://www.x-epic.com"
`pragma protect key_keyowner="x-epic"
`pragma protect key_keyname="rsa-key1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
leVVj9ZLEIHNUV/zgBPPd9mbQvxVvxsDbEr1fVSaQlpdz8acJRTfqXzhnfv89SG0
YM8mAiW5vHIpCI6+qxK/WZQpm4eRDYgFkymGyzoNYy9PzZOisZ/6ll2RjcDYCBJz
Jxgb12/3HYHoK7+p9cp0czKh8qY+8uZObgrvCiOahJwSXxjo1bosA0KWuB97bp2j
RPHoc2nHMleEVyx+wzpOMZBBMvPb7ANIzynmNONf5/xN4Sd6oC58iI2JljOZgG1M
wquLHwFaRb2yX4JbnDYo9wIkdhcC5Z/Lwx7SHqKjqcJ7x8ZbYkPN8fwQujESLLKa
W11BCSxYgGBiCQLmHI9owQ==
`pragma protect key_keyowner="Xilinx"
`pragma protect key_keyname="xilinxt_2019_02"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
AcX3skDaLmwa/Cww1WM/jx0QLkWd/vxd7b/UxtrPU9jDTkjsfskBN3enocvWdUX2
A8WZAfHoPfXNxGmcfWe72Uni3Anyo6fbH8FgiYXXUpOIoH18695hUDt8KjeZ4Lbd
Yb500eQlR70QuvIJRIMHPT1HkaPTzx0XVhYT/903TPCp2iYTLS0voYefnbx49qYe
jSQs00EuvsbxK0pR59BXLZdLHQgq+G3OxLyw+1A1ln4irziOUc8l6GuAE86DoQJe
XgMGXYTacCnkKRolyv+pkQKLQ5UnPr9CTtNtYihIx5hTmGKFhbWNjlno7BhWI8in
KtenTANWdQ0qnafCZBtf6A==
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`pragma protect key_block
VgKmrspuOJuWgfZ+r5vCyOc6bsUGjRW4W+Zm8sloHN//FUvyxVm+fyTkIjleA2mX
nZWemg0OuQ+x/tApRaSKvPLCffRjQs2K3bO6snMxVxKpg3t0Q73FKph26lkpY7tV
r2saI7NFUetwrXxBLUEvQjaozjELDrRdKwhNRzQkJlE=
`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
cGgMbcbgtE+YiqwD3Jx7IO475kOJmKZQU2WVD60dQSpIywFJqSQgHsj9AluXnEol
AQQ5R1is4U9TCRmtcfFLPexa/uP1ANYWxRmCviU1Hi9HKYbhwhusJH2kT4VWDjNw
0XGSkOpH5g7zq90HhjdZVEBD49SyHJC6z+uEETApU/GnukkzKj+Ue4y7XWMXbcer
mprIEybGgDijIyB59/K3Z6mNoNfbWlb0Sfuor1uUpsZJ6v77FzixTFdCCbI0eaB/
IFtMX2PdoJKDkDjFXRAQHWrJM5qJ/Q/qsvKxidpxXJ2uJMi7IQWFysn1Mm7wF4jF
RBianyWjBQ3MdZ8hMXVymg==
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP15_1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
4H70WoFYXpgDeOoJsPX8YQfvzetoodng0+PcvoTVdn0E/sGWptgJ4GxyRN8VIj6N
1Zo5NrASv8i+BXy2NNUKW/wnQGuE8BCDR1pbR/lkVKPEVcnBQFyQoUQJHvQCt+M8
sKs2+jfCvo7Z7+AMxaNzA75++52GM6fgldzFokiDvN6eE5b/O5TGiPUqARXHAbpV
wok/jtQTbvcDi/lm7ELieaoekEnkcoosAxoubSzEFYdGkGfo+J9LT/+cnbnPs5r9
TPOdh03i9G529nZBLfGFt1Sv6RhhQyCNF4ZVaMXfvNSB9NIx6rxg+HPFNde9GgQi
Eym2SMV7D5AEQ+/ShOrOFg==

`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 13456)
`pragma protect data_block
/iW48xkqSYmEIpv6QhO1hO5lGLjYZOgABuECdZCkThKi0m80wKeMYWe+uwD/L/KF
L9uW94pf4LZOc8qx3iaUW2OiX3DqFN03FrTTJGH1++XH3gZnvweFbCe6UoCKeXkV
u3Iibdn0k1Wet2GzSmuYKZiljgG9XF0+hTs7eRDVkSVUG9ly80B+tadKNhwqxdIH
6XoQ7WdNRIHvtvYNSleWGMGEwcpkXJW7HHX7b3rfWdvxzXBpPxShzaJ/kytjp35V
HQhH3FmhyAudL8huDB1X0fAH+Ho3DzXiDYfzsxEI3Xsa1edfvtP4vUSP/d+w/YrD
geNoLoFroY1bQfj8FGrsPXUD2L3Dx3z/qAAhjEM7+/wVFVhGheZuITFrD/6JCFUU
G4b8720BKfnmGYnPksx7ebihMHzyXMy/0QRXRGKo84YOwLzR6QmFEvfZGOOuWeDR
DViqDlEYqYCus2qQJgDY0Uk9zqvjGv+Zwc8YOmcQ1JBnC+KUI8M74Bn/T9lO6/Rq
fGL/0mkk0/RggCUvYwpGJ13ttO6ptlhbsh4cG+NJo9iechh3oQ90D1ccnL99e88n
3XpZyfMMv9P7wJkC4E9OydNJXdOP2Cvm8F921RivI+quL2Babz1BguDUA2BvQrYh
m57dX3buFtfWZtkvGumBjJ5JXC5+HEndFZ1ZGJsYosZIMHvz5sKYxhxtkH1MsVFd
NythqfgBtJtlqP3u7d8vXaQ7f8OSUHUMTp4nWKYFz/nJIX1ZXtqkBJGmXF8Xr7XD
bLIWUfV7/Er4VyfYnrPkIqqCPdIJ8/iobHIWL7h+ONWBaFLF7vygbtsoeeVlSrrw
n7Lfi6f0yME2tWB7r0T/p0q9qDiINtduXZErRRyHJK+FixrHS8Phn0DF+sePd5HZ
DdILqIos63K56PPS0XItVWkmCYFR85dzeIlOl55yf8h1e9Yb07R7EGw3kruytiL+
cG+FfvAuWb0bm5UEUHGBqoDfyC73bChHTgcNLflV3RfB9gvwjrsWL4HiDcAFz/GL
kIEqWsZq96d1ADTi1rDyscPfT5cbGKAo3uoNnt/D8dVDo0enNy55PtwX//HOg4bC
pDNKY1aKzmwbeK0DwtgNIMAD9tu7hXqSjZyLoj1wmcVmAapnk5rFnMuCGTOR4Eal
Yrbx18gVPSlEHN+aSLnPrimrWCzBH1UjyUjQPFBb8szJvBIZewZBdllqQfAYpmgn
/P47VYEr30PvP3hGB0OQ8Nq/o8jykAmRFbvsZhqa84QYxijRWN1+mIUDVEJE9eBp
7BFVFO46tL2tkkLxL35Z2htQStYaje1hnOJHOjs6XiRobdpgjNK6ES0WPsTy+apK
GNLaFrgoagh1y7uElvQLPs+LotUG1HdjwIkxQJp2CXeBkQIOGcwfj6sO5ZXNLdeF
GpUfUEykLL0cL2LGcIPPd27HwDB+BUzbR+nLaxDGPZQ9HOZLUz6MxC1oFFJsahT+
48O/29GdGXMPrsorfnUzNz402k2IrVhlXiHeEsGVcTH0iPkLPM7+5bwsM0mCv+0h
60LAj++7fPLFNDlwUZ+8KRM85zgPUr58vpNih0xgsRKrA0C8llBf2CDI0Hi5LZsS
lssU5p8gO9ikQhDPPS9UNkwcxraiiPpEjv7p3z6gfDVhXezvSPAkVpeZzfBXVqJA
O+tc63myPxwvFGYJn2ieN44IS1g3if/8jrMp8ZUo1mUSUVOrGEeg+P428a+mBWNh
PSvtoLe5BAz6xu3HXad89aTEWCfj7dLLKl3hslZmI+8ldAbKiQfTFE8Z95GVK3lL
nQo7Vv4BXfV5QvkUJ58m+c+Macz+YP4IW7XDkDir2D0o8LVkIjNowdtujZFbd/YY
72heyYib42OQfjsPBl/0Rmp6FNK/I1uV3IHUWp1sIdUFk5Dh7Ce/jGH7I67kHbJD
JVf6XwjKIlZ7ftN5mXbKqs2vRBP31rM5JiYWwnXlPbv1MVRi7189xxSrCk0UZd7t
4OU/S7OHn4ihbuAG/fL8QaucRvadqDn2MGhnR7it38A8lmg7MLRGOPnAzJYVs7PF
AuDvVzK6YNeKA/qXEVpstB+kqCX5Ed+sz3y13S8KXPQLt9G8Mn4enhDtGclqvH8s
zRZh+lKdbOWTMPiy8nAL7jTsvgrhTc3FgXZsvl18HnwdyU0PwFDCMp34n1r/A0rv
aOL+KT0PBZxsioLUqFuXu5hScRLhi/FGDeyWWPY0lUOxgM1ZmAtih68cnU5/KDsJ
yE2qU0FrVl0u4OJv3MyJK5h8HLjA7/IwVOB53mH3Ia4fkdweneUvWBHu4n4i9101
PB6J3CuPLrSw+XZ+JqZvf37AE4eS0VsOcsrVS/u7H2FXOQESmR8wtjREAGrnvawn
UmtraHZ8YzCeoiAHCSLUvoUjMoMZZy2l2tQ/kmRIHqg8GImKhEt2wt+yrPcfBjaw
heW8+c97EJ+H/sm09mnW60uI8DhsgRcheOFq9Su5aEmydFzPwMxKcOtOEF+mAQck
X1yPEs0ou9BL4z3enciJTWn6oWcNLY/bMPtaggMf1U0hykgBSufCm7cxJCIiwIRj
0oUZjXrIujItxeEUv8SG7sXD6D8uVcApm1Y3nddDxgdVUTTWV2Y/Gx49foosbJmV
yvnBBsmCYvsxi98mjQGFgy9Azq0JHQmBD7TDpNCb8jVutWyW8MPLWprjkAmL1COB
uDoHnsnCOI3JlIwUD1pwoIlf3ySRlmYUDoZvxK/UMk8AC4qrRfUHbAm0MJNe3dyK
2RM9jis0eVHKthgQJUwpEzoIpmkIiEVm4RY04wK+/ekrqHw8HNIoE7Imo1R8navD
Xrx+aWZUTTLvLzbmOmKEF4RNTzzG+7wOnm68oxqvH12Utub+qVkto6VV3QpnryQ0
CCku4ItsNA1l9VKKqKppvI2Ew/nYYPS5tDV90syYbeuFA8jXkSSK46XMk+t9YPTl
aXbhZLPju0f296TcZ9/bH9zXzEigUu1ulQb8Kkj/Q/n/oD7aKU5DYKQ7C2j9Ymex
z+/b2k8IfCqfW/R6UsgK/afrGvkU+VPbLycrRKxEoBTpqK+OdSixLzaipSYK4BOO
q3dySBfolXVUG/iQCZw3hgw5Lo8QeY/1ol5oB+BiMwrLJ3XCYv6KoMzfcqorSU4x
sO32OHMPRrXxMFHLLC1ATEab5bS8ZjlYgaBZn/Q1/x2vW27sCFqPPiqJ3w/opf03
c/icujSAWR4hua9wPQ0cllBHx6jCOue1kJi//ocgl7CwauEaMlwjEKhJ90NjQ6ib
1tac3ijEjuuoNl34qM+0pC5oQzkdJ8o3N4laOehOTMlQzFQrd6oVFNOqeR4FxsLM
mVg7xsBsd6+GUY78PKqhI1I24DL48Z+dSzjT2cKanW8UvE8+bCmcdoVK0SJtTvh5
vUwEPon1lSBoeKgGyIqLE66hW3Zae1evTcUKXV+dKxe60urfi8P1eJUBvCHF8iIg
QnlntiCiMNVEVQm5kiPvlWIcz/MLIgWB7lzHEmUjt756i+RkWvfPeBXnotQ82Wd1
88N41U9hDe4MyMSWoZga0Bc/s3Eq1Bs+52Spa4HwFHuLA5VupokDOil5ELEQxego
6wgF8XAcwQ8+rKP2EPNzHlVzrkNcvbYdZ2LWpcliLPAQu8MekugmGXXaI7XblOlG
NDtS0zgccY44GaYI85gDDeAlvAsjTvkcVFdJVFk8ti2hUFWNY3WuQJNe1kFNzgdO
1CZL6IDxwDE6kaY9qhdtaX4s82+UNSspZRCNckfKaaP7pSvH88IjDLpe88tY4JwM
MXveFmtKTEu2EzIX0o7RKDU6fOaf0rvIzl4rligUUHYiJ5PP6fmbpIWUlY1taDKc
ifHi8UqGpr2KSzqqZmoXnX6OyfBPXQ7kLs2PZz3T/61+o58EhcnW1L1HXSCiJIiS
HGUsh6QHt/MkjJ24eyCgs/su/QYMzl7jwvxXOUZu7X1EhApGMYEP7YG5cyruhblI
Xsmf8gLcRFoY7vvHaDCEx7TqGTPUc+vBZ4iMz7HDFRR2T5ywgZpuFO+4HUW4aJQt
K7BhdunX367q6SNHC/+sS8NIYyx7in8mZIe8z167zMMGNtSEo34dDc97klf0MpwY
PM5pecEAQqbJHj0DixtabwGyl953LLjG3IlgoaiLff6brR3S8JMmzSVogTjKZY3w
hsuH3YoFvF/TFAbg5IewBnadxljWmdBmcmFNi+HQS9TaxxfY0cG4qN5KcpLnx5ig
mr8LY5nPNVooMbWnlW13sz6DgF07l6BKhhxT1yxwQ7adQLfF+OxtLK/29wqj6HUO
Ldevz/3HkYCAtVL+EG0/eRPoHCKfO8aW4LHq67hirpScCdTYejfLhH6ruUaelpsw
Agq/KJt1DgaV7rEgegvmouCUuvkc9tcU4hcBRXHXNwrOPT44LcETln6lsUN4WnGQ
ltYuZeJLuzShYuNV+qOs34GEM3+Qc2mzCXiLtB2sFU6kfRM9y9Ml/dV+/AQX0C9+
XdHrQdzn5I016aLkcBWFi9WzhOYLZsL0eZ6Jt6gDMjByvtfeSV20lLyJ8ccY7QEg
E6jtX1Ig7QxqD659pOPLQRlyQ02PNPr7D3jjtXTCewRcfoSsu0tanNCpY1rSz+Zf
stGR51D09CXI0Kq4CC4zeRiqIdAgF2lGBexwd7Vzy5JU6JMYN8fne1VN7uI6IcSU
z0qcFxTzgxC9kuB/JY8dIg/jJfDYzXr2Mi1swuArl9aRf1fRJi77xRflVjZl5Wlc
GT5VYkTKVMS67ExbVRudjnSNDxsxbGsyv2A+Wd8w8lBfFy59fLsDrH0lBWlRJzFN
QZyEnsB/pQ1YXXMkwjHTO+WIFeoj39MRR9U8AHtabNTxgDdCsk/1MgP6qWG9pbdG
BLe99SAOVfpSMj+5d0JzEdR0v2upXD+Wp16EfoNDlCGbERR084EC6Iq2gI1yej5X
kX2E5/1u4vZwm1YRZs2zoBv7mfE75twDazmAtuaXX0hdzeoYjphzEhoQaKJ0Tieg
Ya/XQitO1dBYNBO+JBBuUA4pjRNAdsfsFjj4QOp3u/OOpKxYrvPM7k5c6rmdbaHl
e5vXJXDvgMyp9E80oBmKR031wZxazzS+v5BiXntl/Yf3oLfr3J1LmDlw+rwR7HdX
ecyU1oTC2W+RLt47MUz0D/HfVjABxqksaemK2FnUsvQ0ZEAGG8Vj2NVjCMR9vDhA
RRmuy3NYH31vX1feo5wZN0ndWp4T1CqSUnS5qgzQWKVvkLxDGFur03EPtHHrasFe
lIOOz/RE6Xox2z2oGA22m7vtrBMPpLPdry9/Yj4YAum3E/o9zMK40OT4Zy+q/eTw
nWH6IqYSt/omYddalUWGjH/QIu/UKYwUD8vUSyRuzkVdW4t/FpRwzqsk0vxUvdA2
PviCjHLGe6o1ZkKfMZH7lK149SKh9pGcADNolvFZTxw17YO0H6Ovptim926tUrSO
MrrxbbTR7/EUzE6DtQe/7yA7DPalJTr59nwTLLyj15MDO7cDwFk/oGxpB+MuB4x6
N0qc0CUMbuCTQKEYpw5RtPMAZxiLVRgaqPmrtGsITDwxoalH69osqO2c+bWz6KlC
xpl2G2LvWzbB94TKLffZ6g5AoR/AnFSDIUKpK8kvZ+I4kU4W6dJ0l/5Y8SWdDcOI
XnngVSKAv9c1zj3rY0YOZthhwQPzY7Q61LlUHQxM1JxKA2yInJuhV9+yAIN1UWP+
lgUenpA5o3Pha7xMYZIt7K6rhCSgiYritHmQYQk4HNEgGXWRIMxzMksYhjgQw+X2
QhPHxUGGW/ZFjwkq1+4srX7qOauaHFCXG4gRw4EVo69BD4FCAQy4vVIJ/1hFtOAD
uGegOgncotKt1lN2vrkkHEC6lO/JmyOT2xEBL6W20BEp91NqHmm6QGVHGtRBXqd9
TOn8Bphnx5FjKHVZ8Wshj8u9fcNOLus7IUJVLIajR+Dk4fJ7cPH58N7aM5vz/6aH
8kkV7D+4L1KvJPQ/++qVWIlmuFJY7eqyXxiS2fMCd8dQ1KVf+PiCzh2OL7CYmzP8
YIxICICIgwPb12J33ESWHBinq48QLu53+2Oz1Uujyw7QwvaBoLcxZLcyxzbkPMHx
FrQAIVng5h3htUv+TCeqBn7OYZECXUBIbNuXCQ0vG5mZYNBMkMzAnbT7lJECeLnj
fUYnd3Y6tamFA1X8AT9V4HWjy1LjbEzM7chl99RHJc5FAGM7ifbjA5naJahS0GW6
7wOigisZeqZQntM+ie//h1cj+39JxhD4Y75+BDr1TUqF1sUAYenFUhHS6Gpk9jcv
kG8gcRk3EU9q5lcdtF5f8NwYpM7YJ26ptfB3HdJI8xv/hmbWWDuFsT9JycFJMN49
Dr27NrkRhz91QWdtbDdgkWrdX0EQDKypUb47Vhl1rJYfBAx8BjS5R5EmPU6bLt6o
4aAIOGDGnHCLbJbZOmOLWddkWUxiuCHpQPJEed6l1pV26Y+SSD3ekXs3Rt6DOI+x
5NDuPzyUeqRvHEfJgWxIE+l9wSA9OEqfFi7mCinxgtFoK+6TYAXXL6CfQmKC/6XN
88owXFvOnP8Klhm7sx696fcNaPw8cumJtVfnfDZbYPPxkm/xiWR4xrJo65meHRz5
3YlHcRNGE+MrAREFScFIk67lnTKmuKK2jhjldpBX0YEQnVro5kyI7YCkTjchC7op
jAAAEhxmdt6nrg0HzcWx+wTHPH8eB57lYPaCXCiHpcVWs8z8BWxRzvifOJk15AgK
nmxRoW2/njrh1BailXun0b5U8fozTPFdR89dh6wqL3Fb37lwrMI9pu56o0V9bWo6
YTvY9XQqwXv3R+MLdpT90mMWR8tfR+9ABm2BjqJsXGzVGVBaovYUQWvTDSyOmBii
kVGSNEwdJDPS313ad6k4yeZFBWrQpA9/shLKbC5ORvQ3JUc8243jBmW2mnJRv9N2
iZBTm3kpIZFJnujigjg2hjMJCel2W2tRK8oSBme9jStdg6crvjyFDnNsEePVO9j2
Z96TNzNLttk3ta90L3YZTuHtoZ/di9gKe1+PWu97iX+5iaxF9Df+20MtNlT2JJAT
PbjQDQ4UyK4QvAuPgWPjAp2ehqC2M4gFCttsT5WmbaBjxr1HWSMJvMt4uTpbNctF
nhJGY/pN8IqTMyvcOE9jSiuhSndPcJ7HJQElEQ1Atzy7Uc0Pn9l4I6UEjEZDlMQc
uJUtzDs1rRU+m3qdjwLPoB0FtmNajcJguaWhOuaKw4RqeWqqYsbc7pm3d1GdVrhL
P8UGkm+9fp2scwpZ3UdLYE/1VRd8jnQEqhelF9Rro/gvN9ZNcEkJVMyt1HnGrJqQ
smwlJSDeQQOWSKbhFUmA9Ii1n5CANhNSV6kxigHzkzge8GekHyjW7GhwOWCvFPCP
4e4jpGGKiLPgsYM9AyPeVoyphUp1JPb8wW70wR8dW4cAHkEV0jPEAF4LjvL0e9i6
3F6h3RDnAZ4bhKKPyhXIdhPcSrvOTw8NVFyeu+8vzYu2kAHk1e+eK5dhbR1vGIJa
fqYe08G0qnFCfGIYVJSvTQGhqXT+bq68FWndNYImikkSgcDirkQcHQEzSKx4H5QX
8clxP7j/i/ZRfgjRB8HK2Q0/BWId4RJqlM3FNCHmBRpUDuS5/NcavHThXmHGogPZ
lSBvJWjJxlFn4laoo1XMP/DDqtpS9Ff+evclvgQS6J8Xhn1z95vSauIqKnm/XozN
eMK5V0+uHHVW69Kh0QlGNdlb978X2HmqYe+XUnBrsP+tYFGS6I4hJ6w6MUJozjDE
3TXdU5282UTl+Sd1pCTfOMU2XsXKB5CP2v6NtIQKJCwPaa4eh+60opq/BnAB6ziD
TlPzYlALjU/0FXIqUj32dcd+zT03szWsFr9jZx6lYSqaVud5G5q+2+/EK+BMLPs7
Ml1zzVtnUaUO/bkoLgF4D2W/zCuX4fDAggg98SXp/g9X4JqxjfZrscRyubG1S288
1ZbRljTWoETOW3zJI5sPyMeIRgRCuVAso5fM9GeepN2+bD76ibEqV0HFh069DRwI
Ki+0Z0Ti1tDHvtL8Z29na91345fYCNil6choBggxrucG44IJIUVZPaLYQYhgRSoc
M1lj6HI6DH2z7RJUAlZZstNKTasCuli7kPKPXML9bzOA2cUa3V4JUa9SsAyrNHNH
63isK4cRotky8I5jjAcdZVJIHXcFB0AAD5yqf888CaLrBs6TJ6M5VD4i3+JzU6SX
kRvJVNR+S8xcwEXlC+inPAp6T2VbNRWMFLsx6OOqyTxWtkJQK3Z/hPvfjZ4t5c8L
TSj/ZcICOBd8NEJXWXQqRuXG+pyuMbsLYosK8B5YTFzXQHVU5552uAqZXtkm+MOe
V/L1LsUXknmgB+OlIHXE75IkdQAFb+hr5Fv6Ky6zCzfScstIo++wd+x7Zdctvykf
Zt2X+RbQZRj6hLtv4mjAbs5bdSgWwxKYhfoh/sFcEM532FY5LIVEQG5IrTA07Jv4
kctjjnKQSFuHNK/x4xcFIbHYeeq5CNIx/dCCUXunMVShQEsPZl4LSe/NrZ0wk2Q0
2Ow7TZ4112QMVr1UinZvN392JpRwElUIfdRJ88t3K1p4VIQ/+s6YlrT5reR6GQBb
u7aRJ5zWT3yjWjKLuzEKJ/BMbUu/+8IJvwMutcBdTjbZaw3tyUgzyeJ5YprZM0KO
wXh/U5wmP7IZp9SdG5vZXFAgT3I3/xiTsngQmyJ6lWMrioOPeVUhWq+Ua4SFAjY9
E7H544RVDtZknlkUSUZ28PQQizRnzO0FNBeSOAXFRYgn6V2Luq5BY9LGxs58TfOV
Apy1l7v7y7ZTxrdsG5m/oCfIjRhjEaJWX4IT+mrDE/kyadaCg9+MZ7A3h8S2pbj4
SGofwn2wThCwwpxrCapJK4GoxbYgZ8sTuhdLa61Cbp0u+9uasYvwN5CjXGem272S
Khx28ar4jdrHYhhx7ydBsMBWzpvYrKbpp/Fmtm2Gf/GsNargmTZuzTYZ5Tl5/o41
q7T23JezT2TxaPhtDjAlxDE+ekbEVXmGrzBgTKpghsgqp6MZ/NLYDnpPaBIiSK5X
zrs/M391DtjXZ0eiUJ+PJyay6lRUGKjbAcQnYpHmGeKeY1p/5aVuwj8M0sArt7M8
x20jHkp7psNB2Sv5eVsO82c1XQXe9zBaeFO4/W5W0tbhqjZJfpKUwkO+aX8W+vL0
1OkFBslad7lD4E3PXd3BGGjS9cwnKoVzgqGB4dVO34q07I4h/zJZHK950s6rFUbq
6Iy0yEBqFbM1xZVc8TFM2/ZwMTJz5n7MKIgCvcmyJ6lbUS75sBVGLQc7B2PuHQIW
NfbGHjJvq5PbSJ6nQqOu6cW2dUFIN9m6Rc0dGPJxCdws/KTx30I+jTQi6Rh/ER+j
b0eGwTrZaidjV22jxBlOyoPTmLJWTssMeCmxktiAjhAx+vT61T5AjaESD9KcHCcB
AWL6WGkzCS8XcxHe7/mT0GhjX+YAR8sX2dPpKCo7xdEg/aQOpGwTsID+8eCjUpC3
RGpQRxbPmp/p2SBgFAmbX7RZtLIo5qKYrTkdRI/VP9bA4RQjmPPwluchUblnv02R
93Xe6Om+kznm7HY5fLLVFp39exMhVYN/2785FN2y/443ZRjdbZiRgMQNng97UanZ
LxQP+bDxBnum+DxwOMSvDhXV8Osp2aITk1GeqJ9iiRrts0dCnZKZpqa2QaLF9AuE
BsIxpdeBg8ky/7MVhybQ7ueUPxampHUZJ/g/dTkt/Cy3f/jfdj5Nnsk6h2dLRgDt
78BZmHyhGERp4HHhnU6ZHJ9brwo75RTJPeu1W/g0Cnvoo5nqZP9VH8SexxTAfzp3
w/X5kJWEIxP0WgItp+7jJY1L/6P9rTUT0FerCKmG6mQfh5VNCxqXsFugsYB003IS
v6SbV7Iz0ucshshbygLKnIqJgvP3lVokZOikuykg8R1NGW/ynzaYpwoPunyIHYEP
aFzyX2TCqbgk4XH4hQx3Nkimgzl/SprhwCVhaCQ9qlvinn4xgmzdtKOcoZBYobCu
UesrXETIxf3iWEYcst5fbJWDSwgZkKonsCnBi05O4Qj8o+eW/TglH9Sd6st7WOwr
OYNE8/Z06i+snRk7hC2tv5PKNx0JlI/d7XEyQ7fY0OgfENEJNYlarA4xh7Ibd15Z
mVZ7pWyqFBwjw5JwvWFvM45J3/H9ttezgW4AoYr8xI6QaN51d7R+FjIVlXOdlG8Z
afx/nP+VifibDSlX9OCpVcXglzYuzz0n5F3j3jQ2f/AJL0ZO5GASPBBCsT+nshmk
lkiLUMgjna3uWV6dF0ZZHPIQAaHRJL81k+PKsr1Bw3koWnxohdlErk6rPOZP/RP6
nI8k7OST4s6fY3SMmRG0trnXgjy3fj7KO4V5McDS+x9d80L4dakf3EfsLHqbPDEt
CTUyRfK0qSOZdhSZBZKBksjjRr66n9DxJVQswR55H6VJ5YUNQDa0LsrxBUesdJNO
OKhstVtCIbcpNUqyRUSFJzNN+dBCke8pXIn3jcsR4DNVPba82Lt7cCGrtR2r4nUw
rpyrifE5Dmql9DfZ2UG37Yi54JHXi5W0GFQ4W2UffAa2ed5+dkIbdKDWICYjfwPL
UzukX8iWHf2SfZinlqdNXjBLUSM4JTM2PCHy6xRulhCH4InT+JiTvRWtB4ystthD
za2PquHFpKiK6hG/Z7Jn2TipApLbjQkvhIjw12nFJbhF3ORy9X1gv67Kn8Dv5lD6
Px+NTiTxq6lPH0RvG1GRKlcAYndZAJzSpijErdraXsui7stSGFKV462YSBRKVsjG
/SzUxdYhswGfcPD0AxwvNGNlAj7H31zFbR3EEejI4yxxZh1Wvtqr/t5mezzKzV9/
oFtpHkDWckygyyMRUQkviq+38qgn5I07agb6wpZtaZSdYAzZS5T47yhRv9Yj4gvu
ymdj3W1FkPReMktichNXeTzrsnnGBl+XDRKoh2GvVDWrW8kya7T+rS02p/PGxxTc
g+0nzIcgOPPCYeitXR+wW7/3sBTf3UzHHAB162mRqd2HPn0HDYj8XHRIW48h44cv
CTCsOlMncBf5oDeN60o+dS7dQuFf1LegwH0UnU8oZw89GSa4N8o4U8E6TaCGZmah
LWEk4VfsMIqLmDQK3wXL/0pSuy2O4tvkotW1CKSKmABcUkfaocZRMBfO03MXiDQ+
ty4Fc2gL1pMIT+r+GEjGbl+PRX1+YKOw91Y5lrhhV10Ur8DJqHw5xu7Z1w+brflc
n6bbVIYFhuidnFT3UneDovkaiV+tdZWfMV6vnigKwWKsuDscWnCPpx4xrZ3iDAew
19W3H2MhNisfDC1+FZpPWil8TcQ3LLAI+bt9U3HDm93pwq6zrB9nY6yJVFOqSuJw
96aX8TUjIVFh1yTJnL5dFA07f+O5HT16C1pVXQap+tQz+tGTdwR6ZjOS6eu/ey4k
UydQWzL9WnSk54VETeH/XTD8KkmgsAKeQEyrtz7Wy/Qmx8kLLA/Me1vmEbdgabO3
xdt8a6E8EFlQKs2pHVPs3thVnAWxNs/o5s26iJuSMa11wqqf3hY2SK3J4P1bPCEK
bgffK7Hfa40BDYqkkzby2wuf/xlHgczfqwVCj+I4hrgr/wocjeowR7lu/a73cJEO
E7QDjWoiiHO53nU5S533STpTMi4ylCl+ajrqjYXjriYYr8fqqA/IWjcvO8uGCI4n
kdu5sa8qGDLqKPkB4z36TpLp5xofoalPTgTW0iG2PmjYeWhPGsvZQGqHfdUQ2kQJ
GOr2+LkmQSZnBgBBByTDHYAeb6rJR7QStUbAf6JMe+yrg1QkiDLi/Gxt3brsnYZM
9A61kmVPVO3ck4xBVAI5rblK0oZioEt2FxYgMoTmlZR8GUDAjHI0lZUcLD7oit9E
XkRbKkLowLdZwZ+v+paoXkYyfLG85xRSwXsOKUIuZdCweEy/Js5cJSjcYt5Mvwid
rGBYsf26QGKInGv0ravou6Kxyx9X3IGpnS3TX51JGZrxlIlJ1cqvAE/NLGe1+pJq
4ThQEoLHjsruAOxVteQ5vliN+XWO/vPB+7sz9DBTQGVOEm73I57dTF/TehbG5TrZ
jJjqyZtBNm3iJXqC+Vc3s0vbGpwv3pSA5S4p/tacQTacaMpu9coh5bwsiOI0fU49
AqyB/EQsERpJ4fr+gOb+etj2zS9TI+LySzw+CC2Lyyp3Y1ifhVoLBosyERgyAfgo
vmimileXlJv3a2Ajfnanwyr5teEGarNafFBWnPyEdddzDhsg527MQ5T+0c1IntbU
LExA6QBjmJ9fLV7YrL+a/NldJ5AjdADvIW85NiV6gfF21eIi1OazM29REXdOrhB/
mu8sihr6+HC7LQ1shfTHnFin909kJk4X57mjuQ6H7fikM94b6CRhTgIAMOUiEHJ9
RQ3SmPfHkJbMx3iXQHZ3+PWuICBfhnyCUcyDjP1DsLdafabA95/whB9xPaj5KgnM
YF7whEEVfGuILV0r6qQJ2a0O1IoMPOB5aQgZPxz0pYoH3AG+V6q9Yuf/dkVBkm0T
kG9kMcaPJVemmoGKslIo1Jo+dI89Rsgt1ClQOJfn/lCjEUr0GDZi5W1lM6nHoNqh
jdHEBO610XDnZUicDumJ/T7AJ7cHau4ZgV3eqxOsboStLFm2yoL9dLqjGzTyIUWs
CN/naQH5qP0PTgpWKHjptjPPDVBSYy3NdsgJT1ofxrA/3RQW6CN3nPszbH2+yRrN
48wtA9WC8YeBgrAiHvrJnXUkfTw0Owaxyq7H9WH6rD84JNGi9Vv5Yp5T11lqpSzH
hr0xa7SzZOYrq+ipGQxsKJ94Oe8yf39ru4u8t6i8V5vdHPuxjOnAT3k8/kJn8fPz
ChYdZPxpdmqhd/1UlKlZpUNJNbwdlpTDa/EUkpyeDaknGJpJpqSoR29ZLjXN2lFS
oPHzjcl/2Aovg7S0ZvWCYO7CsoR8Fk0h+pFjR6bGb+Ll+tm+M1FazQvDbKBpaXue
tOMIxy1iQ4e3nNJ2T9Hsc/Kt9Ppa7BJy50YEX3R/O30BMLvGOc5mDiDrKuhSTe3l
ihlWmeutVfH+KHrYU/g6wrgJZnBffcndlx6cMHdK0bpN7Ub1+k+aNgp7tNZIAK/v
6xdgrnaROr+EicWLXXP/2Xx2WT4tAMUcffqhNEMCbhKZA9oiom64Sp3YgjHqMGTO
nzL8KBxbxDHzuYqpcFp5YeihqoSTop0b4VcpzQNIutPSFhqROQo7XlQyqcw/+AK0
x/+L6jKF14UJcgy06zv3ZS88H9/bKhTTHCScB7o8jnYA2qGpGwE/3CqdBdgyZ8Cc
HUUtCnAa9oBHIw6HyHNCcSGvE9vbjjtU0aD9xH1MzGfOKDslqnsp7GotJQUae1PW
kgom87t6oqXudnSk14mblEkW+vItzuHHSqsdqCxeCiLj67cpdgocMe6OdHpuHyxG
l2JcXYBD+ggLwoFer4ARwOyoa18Au6rT3RFVj9XT/PNWzkFPKlb5LsE6bjqFDDh0
s1DCptCHvnDnbmNsoRXOtweMvY2vPMzidij5zzfPK2P6bup78w8taluuJarXMlg4
v22CFU2UCEiyG4HcYGKcYft6WVRT9dbDAc36kFEiXbim1Ud7dN8j4AjIP4kfsCFH
KZcOb3mxL83hdtaXhbwDLTqAU/uFnEVPGOFj43dRFj0tcbS9APQjjwrH89+AwskC
B9Apz7bAkVfSemuM7GMDnv1PrCb26+/4qa0pk35+UVMNGwgefEJ0A0qaYwy0znmG
M/ltNF38YCWZlUY+RHNMCHywE0asFX603aLOhsEk+obQH0tTt4LlVlb4UtYkNX2s
eg1uZFsheXC1ldsrdfP1QpIrqftmol6/oti8o8QFcvki5f+wxd4NuD0TuXw6ST0+
d3svcdh7J1bVaUAYXP8ULypfCWvWlnhNj9DsHvZBQxEtF/W+OBtKomsZT2vel+lk
ezQMF1bo3lFHdZ2p7Hfl5ywuJwysZZCu7v1CK0ouUH75+EEa9hF5BZSC66h7fwoz
RPcCl/rqX9pP6OjyvkTY3s4mA5qgH7egDhNsXlY7mUTVBpEgzFfxX2BVyvIXA+9x
JiizDrCIiSWlJ1nyViNVB964lieR8JJXAuW6pYvwT4EXo2s+qzT5w7CuRCpLoToK
c0cTC+oT6ssVnymCTgJKalIgL8vZ6DBOKh6ToRK3yPxXJeLyrgj5RMCDN9N8xVFz
6qoAi4jKD1rJvO6XmSpzYWNnFJ5l1c8ygX+m04/q3Js+JkNavucIq2Bn4hxH70Oh
VL/BSq2Y+mass86g4smsu4sDvuyPfz2+lIKj7YSYIVlH042OXaWUhoAfAXxxh54V
mSWv7fdsUAE7/8g9kGznFq+quwFzUAVpg6KT6JdP4hxHM0oOkrTxTBnWC/3RRQ/g
FBjaGjdgKKjRWH7nbDqeIQC5q7i5PzFfmCtgXMj8Bkyn9eatdGZs8yaeqvDD2XpF
nLFgjHhv/35/q5yKusvC2rg4f+TkA2wjHyAi2L84eMVQLQkzSBvcUpDa6Iu3V+fp
k1idvf+xuJnKBRiX2iTIwUf6BwzSYJ1NYYJWJ/lcx3xglmJh0/JnFHOHdwlRrQEy
SiNgW1PHrwquu2Zu5nTou/rxHDfttSZJu+7IQUTf7expF7TAxtBwYkRTSEf0l3mN
EbrMn9P4OITaC1qGxc5ntIjEyR1RY+ZUV7jaVwhxk5CcX80Gtz6xQ3cEh+ndMlRZ
4FJMegj92R3ki+BEQIbAYT7dgqFjdXCKo7Ot8fm4o0t0ML6B5pXsK0odXCoLkxyh
ULUkBlHJXnBFxDknp5tg3ozCaD6mmeIM2nGeBmv7JWB9EtFpjVJ3WaSb9GXWnnSs
J97v+mOQ1q4eD7tZtqUnFf/OZe2QL9TznJ2v5cbE8I7u4PhYdFF4TMFei2p9sOMA
18/lfAmMDOjDfxBYuDU8Wzj62CmFPsgOfDlauPLwmZgGjL8qjfKPne5kAaGCV5DC
LtB4ejQ3F9y0vXZtS6UQRq540IsuovOfKmmVWp+12CrZqwzz9csvSbaFZSrRcFSv
the9VlxDxAWqjcu0mbOQMOyVkTLE0H7BTxfaro0AJGBTitI44ksutSioa2KntoJB
//sR2Uja8PR6h1nKsgN35zSJHSdg0/c5xeI8TPrCsCkyUe2Fe88R1HDGXssKGw99
eSs06Q34dtBO+ZCHh6zopJKTIUHhQb+UIJSIszQbzZEuzRSn5cPhjnukKX5WLH4o
P0kiaZux+nWGPoK7GnTSedk2kMYxT1JqSOXs1jrTHLiTQmM04NvkJvo18lhIWb5R
ZjEsqC3wsz83jdMKTWD1vUyxBtLGwY6snuosvTEf0yDwVLIXtEJKRDmy+43yEXpm
4jsu00QVQEa0BibNwy6FR6PX91VPg2TQyCk/37quYf6yZR0tN0JlQOjgviYOatk5
rwu4PNpu4MxiQB3X67UQL2kfPsxVRYdyLb/nCfXvKHIKvi9XKJegC0Py07JqwG0u
dSrB+bsWX/BppwjTTVOEWjdjp/bdmizN4pbdXR+v6Pshe+ll3vFpl7UuK6nz7HHW
HQ3D6M8lZ8M1Q75GNu69WQtEelTtVefCe4WRxolSd25AAFe4lb2NX2FpiLFmrM4i
AVTsRXSVFiw6cNh/VnVMgLo8HGTtcJc6TWSQSLCAmmihIPCiSEEnMM4JQANI9983
+38GPGp2s2R95WRTPhTgA4/yJ+F1Q8MyUC95MJsRJ2EF7V4LQv9Rg9t/7ggSgX2l
nPD+GfuyiiVSY1hEPHlTRSk/Sck3JT2TbzC6O3zm/bxJMVI6WHVDH2JFizVh7/I8
HH58v6YxQDsPTlNpKHGmT+K8Xo3HN92waEA83zSJyp3Y+4DpNKhJeWXswudoY5LP
krKvTyZ5lo/jx22veYNkGBzcqGzzL7j72PYXv8Sez/tzSxKpZM+DPBSotcUFep/5
OXmokfeXGNbV1e3BtLugLQ4HXgJSGG4r5TJR1CJhx6Zli+h8BhmD5O5b3azjuU1X
vCv2wOjxxf96xPXrvpVLBDx1fBcx+5/Is7X6qAe5fhZaaEo9XKlMzGcOOip4Nw5x
/Cytao6/WUvPiEYZv9KHmTZEBszwdgfuNYRqkm5VINg4r/hJ/dygLti940ykg1PD
3tICoYbqMFSkV3MMpKY8331E8NxdHTrIs0JCy/0bXDXrz5fESVMab6zbfACuLkpP
aGVJ74o2w3vDX/o+QGc5BX8C0d/x2dtBUk1Z7vYxbmb2r66Wf9UJB5Kx0OXHVQPK
VNCLvAk3ynbiXRByB37YPCP0+rW1bjOTvGMNivlF1vik8BW/D/5eDfmGfWa63y11
WZ6UysBXnSRWV3qa3yU448AKwhNmqGkCztpUPWhIHo0ECsCSdOThn/SYl/oH07uC
6yY8qwoTiVmKc6GVd2O5ul0TJQPw8jDbNJa/EdYvIZi1kC5LC3CF8YTPKNEKfNw7
qhlzAos6nbcU2S+88QGiRT5X61/F/4LD3Htk36TGsep59XpFiWUJQW+GyhakPflX
bxcVjfhnKOjpeZc+Zh0Y2kwL2b9rtoL91kTucX/9ntAkxYKRcqWNHp8D0ctkYqJy
zZCVk8xjqdkNnZJdQ+sCvCnf5yWLIjEYwxMg4K71v1oqVJpATVjVV4S4LMnyGd5p
TtkikZMKDC6sncDnQv/vnjppOc7sia8hUnMUk1CGzKa+2b6ou/LhKppkN7xzTwiy
mCSJgl7LtWxvbupx66YDoDWJDi0j2E/5ctUhY4M7aDjzu4lM1+Y+2J2HcKZptSyG
z5TyVfvY9WsgYUTQh8w87dUCnzOi27WJbXom+BG2b0RhSbNmW+QcgVlMF1qqBWKB
nhZmDGvz4mWhw8goHkVxSqX6+WE+Pnuo8OkyVlL2O6s2YfleBJpmH6khDtUnWa7s
uvUiEWQCCr2wpkgiwSxHznwl+4pZ6HB2rcdRfRrWF5MVto7pYPzr+0R1UREyZsv5
XPl/PVMYBzsKLJdu+rzkiMBt6LlEypqrFDMfOA8QTtwhIefy0SY41W/GyV5AFxuI
YfTI6zV6GgNmCnlxd3Z2uixqQi656l4pS3ppwymJasy/N8pYuWNvhqZRJ0WfffaB
oaa4rox3NrKPEpJ8/IcRgXcYvloId3WVUJhuQAmDgkde5ss5DS9RJklHNjH3KiEa
4o791S7TiwspqHPRZSR57o+z2OxhoNQI76qOYe3fXbpVan9L3WFYuPKlIedtYyyn
xrS5JOsp92B2qWWfu7Hl7pOFuIeZQFWtJPHCX/W/PD2ARilPzFYELSZuffZ1UWtD
4M6reJ0AI8ErZD2eZpu6XHROMSKqr+I2HZ1Fuv4ylVoDnU6XigMb+Hd/i796lZ6s
6BMKS8XxhKd+ZSc5ygrIVSJrj/jHmZ+ccWDD6gQzzbOHXo0rN2lAuT3bUl3TCojb
CXJrlEzZoN5wOEWa8jkpfKtnhFbZ12kX0B0/rHJ2/ukQo2iCBs7BtAwJHeXIYvmi
gd7o0+z9ZextnkT4vfdfTw8AITB9fXSIyA1rzzy5QSIVKH3Ui2YmiKzXpRK53xUh
P/LxMFqJvmvbg3ekm0Vq6sTFDf/WQezno+md+0VUxjk2/X+2iZdZnQq7rVwX6yLa
tUjWAgibmM4eFTiy9KoYUIA9cdMd9nyEULrCAlygXDCfjXoNzVLi7D78bCj7Sul5
9fCRYPGWEgr8yUsOcB12avpDc62I2oTzu+AH1Xf0AZj3xuLj7NAXR1ALh57ce05x
Tf9lkxacvvPPwSzU5mewlQT1y2OLvIjviZaPNS5JrE72/kaU76OlsgSyfk09A0Zi
HOPRuOj2b82L/RQCjVDUW+Jh0Bym6Ab2j6DUN2iRwBnA4PtrfbwJZ6cTLiCvCpkl
wl31x559VqXerfOHuG6WibCjnUBTt6gR7dW4cGWbmJZtsAxkJxRyi677hheTzR3x
UajTi2XoxcSMvz0+IuTqDsDnd63aaQXQ259ppDmUAzeIsbxnmWXoroTp66cWNodV
RBxaEtxwR5QKCLVC5bjhDA==
`pragma protect end_protected
