`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="galaxsim"
`pragma protect encrypt_agent_info="https://www.x-epic.com"
`pragma protect key_keyowner="x-epic"
`pragma protect key_keyname="rsa-key1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
hvXRUcKi6gFE2BveHOfkBJJ0uIad1DEOlqm7Ia4FZ5gpcFYISh6w+9DNdHoxzOFD
1ZK9D3Kjw7423pwWvLyfoSNAwIgFAG4hT7Wm5S8QWjljRPZDDYVNgXdw4/cxM/xD
x9mpuXFCj4W6od2O4cZDaYn/tPnRXsUqAiwU11Og6uPd9Vo1KYt8eOIp1MMdi+8k
+0DzX1EAmoZJQJTgCuy/IGc72+75sazK+GTs5oNhOlV5dteXQYoWZ9agIufzhvdv
jU35wK1yTrImD8/+7fuX6UuImFNJyEFUENHDwWzyPjJ1KS4/6xi6m3hRb86WM8K8
PoWHIExQlHbFiZffMT+Y7g==
`pragma protect key_keyowner="Xilinx"
`pragma protect key_keyname="xilinxt_2019_02"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
SLiNxmawhqF8QdU1UA7Rdm5m5XM4A82/n0PW+mDvE72aCUo7RB4NccasgE1ffztK
PTpdWu4Fq2ZohEKawr8fbShq7lDF9TLCiLnkUWHxDqx5WASyGQfyUPjv5It5yDlg
1XskBRt6Uu1dn8M7xHzXzzvevDJ7OsDkr9puPhDlAHPS6XbyxsiUEUra6dr7RvB3
/3Pnp9JJpMIGkY17bz4ynIeplwL/H9R04YTBPgh9/lD806fUIxMKkGiDaN3f0rx+
6xFoGG36RLOO7hjERKg6Rq2SZtPnd31hFD/jhhdMT2v0rQTANg2L+xFed5jXqvcS
cIvvnhHHo+Ry6yEHoWrI3w==
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`pragma protect key_block
KQW3BG7pk6REVR9RW68HgFCWNkSn0awwNu0jDzbQUmxXmejQiT53JSIqgT7nR0Ci
dUavRgV8ODNwAGS2Mwm5fhvD7Ud/7ZefhkAjcEiOiThqwTiK0mgKCGWacqecjrkX
PZunWr5HvHcPACMMet4GVUGCWtJDg5jHesiUDQIxBko=
`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
S/fxvZgGiqGOC2mfQZXaUjrPUkZfp53+4z/oVeuzqipYodGkaRlrP8PxpSpiBF5Q
tzjDunHpi3pcaAFdNGp0Dk8o1iNxDNO1ttkvf/9ezavr0y4B4rGPIWUcDbgquaoZ
IsYz376RrwbtEb3ujHz8rcbU0pvPOS1CK+/0s4dk9Z4rcTQNawly4cEDeJQ+4R3G
uiJb3Xc7jMDhWBaAO353u466kjjyCLUhW4LT/jSR88puiprykMhlD4VcfvdWKhs/
5U3cE9IOcgOSAlU8ZmESuj5pTXknJ0YHsCep5w9hVbFOAz+TeTi6LRNj5bidCUHM
I2PmtX3DyPu40inFYfPJGg==
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP15_1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
IScC1zKvOK9M7AFQnjg20wK3oI5w2B1kzhp7421M9OWx9XKbcZGLwGWnVcLjcUPA
YK6zL6mUSVXp2F7n9tEevjwkXazJdjKs1virdOqP1L0M7u6MkFMzLa+bal8LVRqy
btO+OHEGR5Y21mxWzQgA7lkhGCpJc0JHyxtHMgeVV7Q4xIUnMByE2XfGXkuV9PEE
VpcCM75/1Dz7EOfmJ1WOG5tAXy1YSoTvG1LsQOLpOumfkvNdEA/afJbdf03oNOIS
styJpjfIeStxYJIzTmlUHMoGzwQ3oiyLsx1Fl7sXZsc+irWqKoQomYZSqOGTvIc5
B/2RKlECUjCtaYC0ZyAWdg==

`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 17392)
`pragma protect data_block
iTWSsvVSX5hL4ts/NstIF8JzR3nw1+blyvY+Ythn98Whhlq5vKka+Z0/RHv/szEM
3v3+33nCKuz2Pk7ArcsiFcmIQCuFX+i0e5Z0vr1TfX+Q2v/4BTrn1bXPaaOZ9LtR
Ev0iknHvoZZoiQR3FepYXJaDq/7uL8HapjH6v4w2K3DeEtYbbakXfazcZkssMgoV
Va4UscMvbeON8+B4+TRW/udxeeev0/viYzwH+C72j9A/TJEfVNDqqhwv6q9dtg9D
grTU1H+rx3KEUPFSuil2tD8SP8qlkZ0Wo95Rz047FJG1ZYsXLjRzOqtyWlX74Z8X
/de+eJNzfeNBEeDWc8F5Fo5i4RsW2vSoQzabEBxtXAHwF1Oq7Nx3cnyB6Q4TM8ij
IgGy0uvxqOG/jO8otOxXOG1vdXgzvo6mE0ztuyr54mzC7m6p5R6God3IVHBQlMuD
EvEICmEQlOivEd1GClrdsJtMbjEHfGjjSxvrldF6evhHCjUuvcIV2DnP1HHgpxQ9
65O4v/aAi6DUfomCq39/fZoVgq1IRImRaAr8x9ksQSF2YHSJfO/h5cHgSN6iJfwv
q0jmR+D0UyNrbUIot5zJVW929DZWK00gwbun4MQXWXX0nILpvrkmRF8+vuTdeLlO
bggniHQYRb9dUUrImNldx6k60qyrqq6ypdll1+fUszTyX89aP9yTb36taXHyMJZI
PeFDqBXejkAd9P4aTapQDIiI83P40oPcD2GHBlJrmpX823PiMPfEohXkD+TxSdB1
lQa3usjaOgBTMf3BD8+NgI6n38cztSwVq75N6sPjXlJwIEVCZDM89s+2O46Lh1TA
gDsUSwd8yOGg1k6qDGHZBqSDX9bi8s8KbIicebTgI9RgWTVLHEzPE/XQbyVOmye8
CnPrCDKu/OgUELPW+6eTdeDkavMkyEAQ59VZ88pon+Zmlgwp35Mgkh7I/jZOnryF
bYPIydu2fRLucpi9H2LTcY//BOKEQsFMY5uDFiSeN1wI+AHriAC42Wsqel3ic7Z6
+NCTYiOU8HbbLHoicjchOgDeo+SMUgymU3R98GEKvDz+gPQYTVgYl1FEQaSx9ilQ
LqZPEVNXaHchN5M5Y/nVsm9ECiI+DKg/cg62DVInbe+orh0XXb9sXTOizOi4F2gq
c2kBf5yg+SxcAp2VoULv2iEXaR4r+o1LpuBIr3iroMVpNzRN3B2nwUsdZcy4F1eA
m67U0PHjXO9YwN+hSyh1Hcg8Mx5F9U2E/Jpe7aqb+nyyS3HPmZACjrFZwoxaUKsL
Yu9D0sIEcbiQWqbJaZ4TSzjuDm7FeWXdAl6ceIqInYlGpePpa3KsrdhGuDyhjF4S
Kmrhj1bUpKk/9PXPv/E91t1mVHSslFTEKLFm+JKPdyp7xp99RGAUgQpPcGuwHEmG
JjtJhZ8tQdRT5Y9SA+ZRiNizzRwNkg4Yo7PWCeAlyKsqAxPWidmBaVkP3y2Mrqaa
u6oUxRywDsRtd0Xgc8770pG1ixWtw8M5oBS1d7U9447T5g7/Dng5w0gClIni/5+1
uP9oI/hKhOAnumZXX8SEpMde3ErTos81LEOE8zFJo+5rQEOupZNhr0uX06DYMBJK
a/QW36Zxwt1AOcWM1dJ33R8ov9gis9d1M2OX9Q4qPMZQcnk7RcuPDa7pKDA1KNFN
6cUsC4hsJ9sLxu7re5o1TdfLD/fzdPoWgpxK3DMJfjdLy5TYdbu/Q7eKAS5F1VYB
V91gDiJVGikfDf9yY5sLQ31BgWTp6YWUezmcploHwLmuW5+IsFOARdAwrLqD36Fb
VKQJNzWEWpFXmi5vsLyNS7VPDCsxm7R2uZ4/dpR1kaTVzVowWA6+7si/BwIEs0JC
vLIRrrh46UHJDb9FMY/SpdDKLT/gm1RuG6w2ZjLDTmLWZ83eQ9zemeks1AL75rxc
paCGLgePxmqp0raD6DCz6J77flGsTCDqToxnkPL+FKPl3m6ZraCZfF0xZG8eNwT+
VvWAMyHNLbRWtUtI2v/imvYShoojyGrA4ROMBUyolu6oh1SJ3Jw4GovA/45UTTnG
XpjK8z9cxPi8+BGgUsrLXruK5M1n9TnY4nsJ1wTWtIvLcHoloR7azjSTpBQTr8cI
siLEXt44vE99YWMU7I3gv2oDtIlUFhou0zV6ioT4VYvVYFWi/6PAga2DhTbx8NXH
x512Ok7igQIDQb19jX2ce/XRS/MbPBFI6ZVGAiIeqHnqLzJPY/qMWnVXgVYY1Ij6
zRzBANEpmFf/xZzfqZ6TxnypmeRwmWtyGZ9NQMvluVw75XJQAKXp1L73SZrVwwss
Gbi5xpaC+2lj5hL6c2EuTgBolYlH/dUlBqRug6V19t2XCjQQg3oDIbR7rI3O1+E7
4ly1lFqbk2rfi/BF1Kx/Fak9mD94zAjKpgQIZTTRulapDQgf55ef5jBmTV9ovF9i
kEKWUqKayjfCJoSQN0bGL56vQyQyVDG9LxCULdXsI3hj1w9WSMt537c015N40iQy
JdPOa6T4ygW85Tcv3o4/yY3l76pVCR04PSmtoqOfPH4KsWYaHu5hXmzD6l86eiZS
BzFgk1fm2IDDlQsAKhHzSFjPHjSnh7WqSUFCWHyqPkoU5BpmXelbQGw3sWJLh2ER
CUm0lHSnA35Djhoymrv0UORNuoiU/4VVbQ4HkL/f1XQIikWGuv3PNOTFgl6P/S9n
I8PBnnUg6F+6GDUScK9oEReF9G7FsCQ1DWFnqlUPTYdSYR2HqONS4mQm2jqKNTvo
NImN0cxeYUfAIFZx22oDlO5F6rmH02foM6mjm0SjIk9JSZxra5hZMYAeaOZfkCKK
rMYI6cW4bx5ovHAIhjTPZc7FbzXgshd5kcli1O4CmLJ32PxSElIimPLSeNZBhxZ+
H6q91hpheBa4LxsTT6d1UxBtKyBx+ci6ERAnljtC4FZzxaSTJE8HMSH4CrlvF8Mh
Pgq565lLv2aeHc0dy5wyhq6fSYgjJZwXZsPrPYxAGWLgs8IHuEPNl7KZcFYMiUdN
ogcMhqf2ZqKZHZeGa+7vUxeT4paiYRGA/FrzZPY3Q8NJZxiLbtWfOMVlxps2KEDg
4cbZMFKrQjc4gZbfYywXtkLDklRKb9dDdAUCsOvoq7K1spfcHwmSZwK7sIEDQEsC
D2BdSL6CN/fmOjUmw5a7ow7z5cBpzopFu2V0kchGnqy0+VdnD740UJmbO4qnqhF4
UuuLDUzKBe+kdq4TbtcpRDNXouErH2PpIg9zX00y3izqJVY4BU3KjUxtU9I6NQNO
ZqHHlXWi4YY6ceyFXMRERDyI8JKXnhC8r6j12uCZzKv7iacRIrNv5mjxoNblwinr
LhG1gPknD+y95v/8iglcOH57wx7sDv9DpqywQMOw4e7HdGTkJ7x0SUhXQpwbKtPm
tKl8nW8IYIs5gE3/z47Cyzum9aTCOTIQk9tR2tdJV3Hn8FLnJ4OV/y8lVJBg3OV9
YLxLOufiKGoDipP6jtXLO41NSDhellNE8PRGYihyqtWxBWhrr+AVv9tNvStrgOTr
QZwbi6Fikhu3LIywnc/A4fR/YM9GfCNUTtYzD/JBr9cIC64fUmRl3iUBh1B50X+w
olvEK8TE8khUWdwI/yLbvbzowALBXOSDeT7eyAPBres4zivPH4i7NdUa0dpUs7Tl
MaOCUntlyY3erpqhj4zELBL9Sp34XFKg6v6e0zsjVuDZAknAMxW/DPaIieJN0VLN
WH9/+br94q9FtGb1tZD90xsXgxnYH9Piftgnl9fllR4d27BFA/yQYVpXaUp+b+5d
p+/4HlkC2Qg83gKAj1sSVmwd4vwCIWX0KyYkk+Ul/4LqmEBS63JkSpUIRadwS3wu
8kD3tfAvkLIVDl5rJhKTX44QZG0RFlu6ld1FA/P5Yi+PYk0roKiTC3oEAL4rhn6v
br6S6+casRI+8scQbthu4d5RnJyYX1FBl2/Om9r1GQB7PDUaf9BWGm0U3SvIg7Zr
ZgmxDeljrPnh3y/aK5WZOcD6UP1sc9ZTv870CihGlBFzWVkfHDrSsBFaG3xFc3jx
dueb3TTm2lO6xjj6eNjlQbJhawpGzI2EQlryukCH7AC9nK9El+eH6aBl1Slr1aYl
ySVBo5Zc8Wt2J2CasSlX4fNBOeOdjSheX6JNGUOnlPfAUwdsGNUW1VrwRvMz3clZ
fib0pT1BbLAPDM3H8jiHDGmn/+lnsqPYVtoNqDsG0JWQ56P1Xrj9AfS6oyRGYNse
H2vG1a1yihSYpYq2AIZ98b7rmRjOR+MY1LIxnABZ5yAgcOAmZ20FZNEAqvkP2gRP
P3e2fR5xVozq0/p8pHaojvYIuDGJFD+iQH4OApbQp23pggxA6mVZ3ZlaajoYx1Yo
ish7plhucSXGlI3QNX+4djCjbIO8jHgeoDFv3BbLnNJMk6nOcUWRaT2XqcA02LQu
l0xOX2oFoWUngdigX+NDef9UQGirtmZ8z4Fb7Z2F3cCig9tmibjAfqhql9MyQPTS
2FAksGU2s7VmGYuUvV2eI+GOwF7/3NUsKapK7s6SGKrTGwmtdA1ZyGTl2/1SORja
7AMkN7ywdGM7bAzR1rWTTWJxffl+3TmX3oKl63xI8tDnqsWpxY8uheaQXqFfX8b+
WZ0jTOEx7P7qoSVqqtqrirLYMHIuekGFjfGPzoVbW5/Xhn7f3C7YI1yTRTF6TGZt
GpU/VVWBgxA78v66Xlw58sN9pj6PVVxWAAREQM3Cj3gYAUrd3mxNrMvFnoh2lnkp
prx/ZPpBhpnEETSB5YjBurxv4ierlzWuQhKshsiy9A6ioqNjqnZdFpotEekBFrtH
A9ADEvvXo2f4E921Ab4MTBbtPaCr9CNQ+bj64woamVuXSoNMDl7ug/IjAOlH6uuC
ir6zp4CV5/jrlZAGgIZLYOj+7nc3BtcZaUcT72fumzFn5V5nHatbnYje/h0w/3NQ
S3vc3ypi9uHIlP/dNr+a1cQL5+z4isYzn7yj5UlM9+WBi1WgFcDpmd2h6sszTGxH
s+m4M6HWNIXVlLbEbxplsdUFQeVZCTELRh24enD4ZFHiKSunXdNPRCER0qFMEOJy
KA4J0iBW9PJiUuSxSmo2uP5I+0FHelPF+0Ll7C+E8UdDKM5KWCwCaRpa57vqCUPz
2SJRcfJWcllxuwaO8nRVI63kHm8oE9/XUNLGm4aQ1lSqzSK023GHsKLViOxizux+
KtcvnQ8Z7Ikw32UYt1SrxIZYo89U3qWFK4y2JEsUb/s3HUg4gc4b7tdex2Bm3Q3G
mSq2ngW9VHN3LItqEqKy32aAQzr8s0aPRCY0YR/l73qjTCIuvwRoNzEKm3pEuF5B
Msxhg0JhfGd3oXjbMldtB3bfbubwfvYDwWjrMExRk+GgWKIJAxLnbdO5EqctaK/H
ak6MBdC3/q+oNoUgPZyXDQo5JnN0rVtr7sD6ltAyJbyosBaerAuvkh3OzZaKVPJ7
Tpw1/F2OdC2ybdo/t4ffQ4lgnNPe/PcsUAe+58XlGyVpaaf5wXTiVAHsdma2H2pN
54aBy9He7f0VQxF3lBWiiQc+sCq+V2ZCWv6Psl28g7rf5ugYEH+Z41T8+DVbkjRj
KpQMDR60JchtP6IP8vVUo8SU6NbyRWjnXLzP80KIArYTOKCZ/o/iuoFoligexH5X
c8kstama5FIQWccbNJ/xMwMsABqQFPtJYHJZWXa7+928JJ+1W9+BNYPKnW7Nrz9p
TqSDe4opE4sytf+DxTGk/eQBGHeA2cRGE994AvUmwZLF3bIImfZoPO2Wg0Ee+RRh
DroDuXmTWf3USi/QjoVNpzBCMgy+jWg/VPn3H5OrwGqfzMlsmwa4YR6SB6/QpGeC
GWf2BkbDyE013vYo/UPCqpPZQGibdvNGyhw1FWvnG7hRDLVUIlSLTbmSqkzSqG/b
a7lzN1yqqvBNnyNxJYff6U62a2YwKauDWW/sqlnMFN4hGLr8ibvsENkVjgYcWrpK
BvFfP2P96HSSd646PjJpF7ZUuluT789GHhStWAjbVS/4LvMMpY3Y05IzzmJAQ4j4
TXtVkZVnuVDAMzm0tvpuKBVbIHOG020IOl1yvKQjWjy2nQnZ/utLZzjdKsPf3fJK
v5dl6pKPi4uu6zl+1+8bMyrP3A/W9S+5cfEFONTJBgRvohDQzoz2Y4MIOoBGZdit
bdOjJxxa8nrh+6NW0ntJHB2M4J3NEVvZAirD/Lc5XZoIjGFi5h9UsoPR8pv4dWvw
iaCE6Q4PdLgo/cgBXP/X/wbFPNJiTF4e+z+FLPt18TfhRXM8lRM7vb1ka9MxEZ/E
znWRCOYb2Y7CfJnpTiIVaLrhMpz+MTqNaro+4o65HVo4ySUcMjxz3ciwHto7REIr
Fy9Hy9FmA8ss2eV+n3VcWvpDNeDWlpYALtTZeiD8ylszG16ItYbZX04308MyFF11
7rlUNa6HrGZQ9I+S3CmcCb2lVwBCc+2K0zGbxm/OGXM6/ezyfHFJ0wX0GqszDd+H
N8WVj9YwiL5ZM8usDdJBKyE+qyhvIIols+G6gOJ7rtUvl2Dm9IKdmV/IErkroD2l
qZu8hfw95QxUlpzmvEf9mbpnutQgdpjyKpjyqfF0Uh5EENurmtPKz6e/S90TKf7v
47spRgI+8mxFIs+LX3k43AuPbK4h3PKpTN4tXneoAWxFPx+5DTYP1k8mt7dJPrJh
Ln5pdV0RdM7ILERKHvVA3PW1v7qQBQiDferrsbv79XqcSo/WuXrDUdbvo2dUxj4Y
EYk0NAS4SyrY7xVApDv8Ml2NrT/wkdAASvo/YJMo29eM/ICfhzllWw+3beyTcZc/
JIBIYSQ+fC29Axc9LXdE3JysirJaa120zi6ydrwpvrIWB/2SQZe2HtcAbIvhAA8t
Q8e3AEa/xd03q34Z22TlgWUmC8xnKEnKKfpad/NOZhdRqJjZfSpxycBfvKdGfznK
19zN+GpkkI9u8vlN6+7aYyu0dFnWpSOY8s6RPtaj/f+ee98ACI1w/n1L3YBbB751
3nfSWXx+Mcv5MuncZScpEgZ+pIzeLerrmPCqHd8SLl8kCHc98rpbCe9cnvWes4RS
mQX6YTDvgb8SkbkEl7LPcQf7NcOMSy51uMEUef2aGRKUsD56V4bqMKhbAwuOnF+3
W09/DtTq/hEOcTLYMDv2iKJXvaaJpLkfyBI9cepevhkqjQFVgQehvKKGIYZuTiFe
sHynGHre4ZxWTjuiCeGEcBACmWqZTM2sq8vA2bvk0I40eQFjbGj9qgSrElIEr3n9
sejYDSUaAcCyjeivV9IemStS8/2LxqMupd07xTnfCkB3IuII6kvYpjsxTsTUib+L
4oXUo6F2dw1e0rQjpompryVYPnmieMszIhigOSBcvRYF3FqpluxZH2fGBiibmt4G
0N8f9+h/8fnm0JVdiRpDQQW1bMCKWlaRll0ggH8HqMP02Vr5fNNMmOYkFGYA5CG3
wHPvDFST0Y/ZBe+agoeqjNoBbK0xvS8IHatnQsmxijU5bz0qQESCQ0rwNS2NivEB
3kPSNOFwBUFKwUL5mL1G9k8j2t94WBiqOehbMEq1sgfotZ9Wf8a3h8KlaS0gJ4XQ
q83k5gCiCOzA3D9eXIiF+unEA5m92t4ES72OLWdCQVgnTCY8xIjPpB5LolIzbzbp
N3BTIyO7kKt6RCJ4CMG7Otb/MIkGwwZj2CL78Aj0f5PLujPMvGmz1Fj2a2lZ3r9L
mdS6ETG8POlupLAIQBRh9cTgfD0PYNRwoMy07DO+bNQuU+9OaZ7vGA53kgWFq7a/
JH13LcGEQqCn01FbGP8H0iqr5YEM2HEzWuOSYS433n5arpEEgSnTcsKV6T8gQc/b
XtBxL5/ZEyCbcKnaGQVfDDrQErbTr20SI9EXjf1ST4lUwMkmVL1OHoR/DXHMLpCT
B/NQsZamUpZBwqpX26lxyl0WvCqzE8sSwm5rLZJ6c7VH7pFTR0ihyTW4Xqcz19K6
atmNqHkP2MuXeOGa/PCzJbYgxlD/t++slxwC2OmZ9SxYq93V25OSpSNDMz3kuA4l
C3P7xfgIlJrC2dLcHuD6NVmDvIeoA4VKw8O+De5nQGthcXSSB9w9BTHv9rD5knmQ
THXXBYED7CB8ylCtyXDSwSIh1CQ1BS39XjMi5n3mXQCKNJ2dfN9Xf8like7H0ZLh
KGvIYRJFC26+5iDcv1ejA0cjrD1exWzNKH3tAc9/3198CiXqgRXt/cS1EBoOPth+
fQvxLN4McTtLp9fXIwCQUtguIlRP8eAeoNuZGU9KhFrQLSU2W8a82x8spOTS+QOU
4HBzlUSLLwI3Ml6cEjzWZWDwb5KtrQGNSxvBOm4Oa2JsdrqinvAcCnztMrr5zL+q
/hMMZOhE1NQPx3ZdBTkHp6ict7SgPuW6ULbaxmiqB0iP+CNcr/VBvFngjsKxq+qV
BoogVGTs7b6vHqIKiriu4XB6Vi12nFwxiydhJmcgHBg/lBu3gpcefdZ0xX8yS148
c6gHebU5MelDWeoT4g6wwPkSXL+LZ86yNkTWm2zUPCFawQkrB59o7Vmpug74kZyZ
LJYucXZ56NYytOVt+WYz2dvQjHFV1lLwNTU2sKLRXQKJySbvaaMlQ9WnJrYrqtna
3CcIe91evM36pOn+fT3/fOJrlODUh5+sh5ne1BHeNpdjuO11dv4rZlUgKpIXwW5Q
ewNF9UGXvBammJNes9b90ATgHxI1W84qKFtDBqjOy2+n7knPvdfi4i49HSBV+QpC
FRkpSSpN/OPYvg2rP46G8In4cD38ncWyw5K16GAYIeZKNrZpEjK72l5d/1zMx6nf
cw03w1NHlc9CuwR5m0t0C2qGygt5AhxzA3xnhGvsFSSJUgeiTWMyCO0J+8Zd4VOH
CEQNDvHkxY98XPXWdiYXe2j4DeerW+N7XRA0YAtEsmFz4mRvqlBZ+v8QnSOuzAH5
wU8dgaK3P5SeblZPa450BRxBpLkoT9jRV3WCnoZgg2br50mvqMzmyies4PiA7qJZ
ZqjwbmfweXwApSpbeUG+9XMSdto6X47D1ArbiTziZ5Qu6vtv66o086QYP3bSpLEG
nwMe31Sf9scCPYjhyD9AZIUXOYn1WlG04Ohj52H8nFsXQ12RytH+MJ697fFSPrri
tB1jaKuuG9+sCONAL4gG8XkVAaBKft4whbgm2A1bXXs+3tbycKhBwgC2fVAU8lRM
050xdxq2919MlUkt8QDThVcP2uFTwLdtKjpjpJ3nKM4Ysofb7gA1Zk3vWUSEDSLU
S7kmruoFI1xYWSoDUlyk+8aGm/hjRLRuZquu0ieomFzSs+fgqq9Gzk562jIufWHY
04r9r5iIGaaS/vXqpGmtkgI0s7FSifNsvMnp5HswxmwIeHF00xDLrDAstWY9+XIg
20mWSbQhM/HMluhqiLymXpyGdv5hDBDufq4k1rRcjgAFwoUwXKE7HshJbpXBtfq1
8P+8qmJYpDdbeiB1O/KxPYWShulq02JTgDNbp5HNXxxIdWUC7ZLkumPBJWHnhzV5
jfuHzsytipPX6vjs2l/1Fr4lc85GO98DAgumvrvZ4Qox9fZtVGMk0QYQ2SdXFUt1
GIvye95BW1UnJKflY9MroCVx05aP6wIvOQYObSADhCJXM0maSeo0NP5nl/Cdf+TE
IQdhBE5Mbmms6TZxweEkmF8WJ7+cm4Dh9r5iqgDZUAbxeP28h4ZKxr6NZ9aUP+dY
zCOuB31APTz7SmHWhmuZ2y4vFuumP+Ydqc0seZ4nGsowxtGflnseaxLgkXeEdUzZ
ESJh4osw9j47CtJ4zJHKasqASZbDF/PrXTg36WMKeiED0yF7QOpF8AumGyF+yz7l
VZeWTlBp9dCUMcObx3Orfm8Wd7gsYx5jUCXAeQy0B/lWYK9XFiJdvfNEjhie07Zi
mc0g7AkON3cXv97ci+sHdsvNHBUejBzNP9gMN8v/fk0xOyyEXuhvsipKI/lKORST
URVz2O3DQNP07YiUhEF6To0fX5VvkrLAsg37dI9X+h+zQPg/2ZUl5RzAp+BYvLlx
udiNPj5iT1J0kxU/hDReWtzNjMxH1qii+vCGwDFoGVaU+nkJrJYsJxfA14Z8YESl
GwqnPgrRLYr2hfkZaZhQGKtwy/tf8D82rPd86Lh1K3gb4Rp/iuTwE11QrxntZQDm
IUEYJedYfhGryijKCn1zDEHIlweIGrQBfBnH40O3odDwkPv7co/3JNepRmi9Shc/
Pv2pnv9LpwSazooliimJFobcvG3CvCQiR7dLao1/NCRfU3lYhzoVpaCqCBFoZfF/
UTGvngktUsvWSTkjmQlJeCgYDWUvtrVdb+ZDkGSaW1HxZbxYvrGg8wiqrKBEy8fx
LYhZchWFuBFPBZuSfAPSzIJ8G5Lo4m5GjXrW1aEt8R6c0SYgPnsx+uXMoCLzfhee
lxmLMNTgIb4DOSKtNA/hAm45UxyX4WWfK3HQxOEsZIW2+YErgvYQdseq9VvGmU5V
ftl2YI1BFl7Xh4TBv6zQ91xYn4xqP6vVZrxxK1XT0NEmaUI08kCT8ULIFHXDuxu+
Qpp+ODoULC6g5iHslX/G5ExvSb6ND8g1N+VDM3B0vErBAiX5xW/Y6or2FvqXcHVS
Gbks/7Frl9mRyGxUFkJ9YtkNNzW5fGXNNvlB0YOZSlsnaaRXHVdiZfe+rGSAm7eI
D79kqL6kt0bbHwCd3Kc08QnYyqKG6m/EDIDKBbFvGsJIJy2AUb8ro6tsIy2jXGt4
gchObXoswPsP+2NthwlL4BsYL4o/l2NzPXMdrOac7+uPwEBM8zmvmx1vKss4w/Rr
4wIeMv2oPRbXWRhT70bg6yXxWRVXaou3KjphOf1X50Q5txLEIL9nJLSmgSDsGE7M
T9xvj/UMtrDACmRpg5dTrC7fM2jOoHMIJ72uLXMvGtpYCHbBtT5ybzEc5T8VwNXS
y3QOF2C5FVfSrsMeeqJ7CpJcScpvpClGMPXnmdW2Z4VmWXGwPrQgIDv/O0ig0oa6
sRY9/JOmAsTa62jkKMvcqYTe4kXcAIridD0bR2/w+zZrmgV1f5rwU5nUYr4g6oII
lk4OYvK5OuXLwutk9WBlfR/mxzmoNDeEcqZSf9MMHJjinSb/Bk/GSWuoOyvp6njx
imXd6+AS6b371yKY0mylduI/kOv+8LPf7q0ndypYudXc1hGAl0lpazXHa15uZFrP
2J//5tTUjMOQV4cYilv0iZqXPnnnmIqHP2uTp1AtsC5P/kPe9rJF/3pcfyFmae59
Sc3qaw3eFLbIl3eRSwhCr6u9UV/iAkM+TraSYfwkVRK/y4igC/5mXado28tPibFG
oLKmR0VjqffGLFeyfKuhr2q/ZDDDOeftpyd44nF1DjyvI+bLykw76q3DR0u8A5+V
P3CC7pH3wEh7nAwhkjARyatsMOWZ2GQlUiklIpv7UAnduvej/NsxgUwh0rcsyprD
IcEZpyCbz/tCHAZyUdK0Lyf8/Ex/5nyC675JnLvG5IeXhZN7NpQI1Rl5iNEKlqMP
iw8/Cu/anWFFMUjQ9U9thIMaD9LYyoRQJKyF5QO+mXTCnrEvEBE3j5gCfGg9/zPI
XRcuyx1pIui6/MDwepeGvRVAcdojBsiQcXvYOqumigFDJqarOPdY56zr8LSk7IHA
6xgHagQ5dCu7Q2l3WAoTGdDcX6g1U6/BNSiNk96NedQck7yMc2R57KdDQXwk/9pt
X94+JqJvrevlvsp8RzJj9ebgXvcYnak243sriFDzgaScyzCeFzNdhseTmzStAm7+
zvdtkX4rz2eYoW50dfLzTL4H0gdiNFlWubsiL7vr2Ry5ZnX8gBX15UexpHaLqhzS
16lsYDnU6w2j+te48Sct9TDxMYubNBd/I53swZnd5gLajOdh5vUsa/gSL6YqyvVQ
0i7GbCu6bo9Eoi32Cm2q23Ys+3fVORZA7BIoqqvqPRF8yg/M9ubZ3G6n0QrmpL7e
TMFApfvp9ZBvp8OFO2nRyq/ClSOwmnKY11QcR1VMakfQCQoTXbf9Ye/RCsAxieHL
GfK72QGtERXdk+ba52MjnZkNaIRxDVdRO40boGoYn3r6CGVNaGvDWxmhOxP2LErx
HYeFUUaaYzJRxsI0aUYfsjUXxD26BFq+WNpK3/sVJSl1OAUBrD0D1SCAKnvyCYYV
E+NCAdmBnu/eO7YIZowESXmOEajliF43/F3RzBLT6/w79STAlbQPCtn5XKrMRST2
wiTCSd0kh5hrZp5Z67PU0wpq7kQ3RmkqsmFOr1Gl/Kx5Yh4FcUxiRVBcYl3xkVDb
c5XXRLMNo6EX7ShVN26YxxYZeXVVw0QE6FxafJOt5idiTMkk0VuP32pTWI6cVbR6
CVlYvp07OlaeWulnP3Sbd2Ln3GoJLTuUlG+Y4SOOfSDtonWQk13p1O7W0HTYpyzS
WDwKhlhMsxGLLBCh8nC4+UpnSY4JBIfuqt+i+wdWbafFqQ9zvCn27oOnIqkxThTB
Jtk2b876o+VbR5xxb4IEsFvbsZOdR9OcB5R2yB7bixGDP0p7ecciDXXBdrBWOHoc
G+b9Utf26SfpNkANiOmZHPfer+9l1mmfGkAQceAuiKRltp9duNkgtlSmqQ0J4m2c
++V/UZrWOdJBBhN9uKy9IgRcgmO7cfuaWUy+ym2UP+dXPvnKFUV6DOFvJi0BYN7m
7z7XnHf5xpHiOyfaSMJvNO4XnPfphTG2hDiI1D1LCMpAPqy5GN7Z7xA94ENqrjZ1
ALhvZmbfz6GnwhTdDvdP/MsQOpNeiciQz4jNzBZZv33Bk4EJQfP2xck1wVcvDbEN
+ELSkPxOxjCdWJnmOS5eVPKc1ljCzWSuMnY4zvzNiqyr+v/I6nbtD9w87rChJHab
Ymob4wMA73xEbe6szjzdqr4PgH1hXclBwdZzMkxsz/jJaZsIt0HvdE7nlNlX+o0A
Yxhu/RHQNEGOMVXrV9y7NntXFipPWsY3ZCdPbQRv2DfSrAhj5pwrCNPJfVi7QWk7
I8zkNOcW7VZ/3XCZeqvVPeWClszI4k/d3RMhI0gn8rr3HI82uK1iOlY3kO6Fg8tY
5RP7ELuj1WqnLTTXkbiFzBNCh0dI3GCmUElE9Of4pouQgijtL22o1IWhNhhSq5iP
skzy6ijf+QUs0sguwkoVPRt6HNtqdGIOA43SamYKdNYMibHbBmZkg4QvgTt1Kx1D
630t9h0Vm9k/s986NKn4pT3HjD0kE6qSddr4p5i0toVtL1o17incZ7MslvTSZvWL
72lWHp/9xKM80w/BHlCcsw83mlkwE2G+k3KKg0/dQzHQp+LdJgR3TaLWh0feLUEk
Ca5Xyk7WepzfFmukeNL5V0WMjRR9frRJ8q/YPArbl683BfS0rtxF+VlJXIHHMxor
ByP9l7T6AUtV5NohaZF5pCN6RVYJ0DwplS6sr//Wkm7ThVKqavz+xgPo3vjpN/On
Eas2+Fv76lTxtJDo9HFXUKhQmNIekPm24ASe0A9o0lz7Xo2dNlQKlQgBaqcq9anX
r+IuWgLCjKI9MJCrTNDYaG6fMIU7UStY53eYtzW5UdW3ISa7dEzPtpns9ub5OZAQ
P2oJYQjO8qBFhSnH3PYlr0wTLw+Y0XxQPJQrxZt8bgoQOgK4xj3QyifllxXeSvIh
Whn4OvP5l6OMHvmGUbs8nYZSzFyHMSGtidKt/clJHaHfxVdZDDdycKcnCY4u2e7r
LLUqeNvU0QBkVaE8mSCY5nxiOdVZo/AvugraxPhaoMu6bF/Sg9EfAKPCEf8qavQf
ZF6NDlBYE/NYyC+X0/soPzikfxxCWOWfO2jn1kLi53kjaR2WqaAFccGbxPM7ri46
40An0e3WNnwUAMLc9uQ8YHvPG9H89jANEcEc80xyF23nNIkBrid1bdoZ1jiWXUlc
wkmKFdVmGdhqNTzSF3mmEUtNUKNlLqo8Ip35Uewux5SCQm3hhIEcGT9HcqWWcDcr
9bO66FPwzFtK0q4O+9nSRJcYLpFqtnN0i6Uts9nyijGevAQv2LgpFW1P95BwAIEX
3dXr27ePx1k4TKxtGUOOzfVmDJgSYsd2iqoX+LoVYRQAzOj/ojo0U11DiG9hMqwc
/I3IdDaT3e8hB4NRKY6LpdCUEYWpMSxPaW727mgwkgzKzw2Dw4T42C7vTbYh2xT2
t5oTjd20izsrHw2Vb0DzwYOZmrXHDBXC3Dj/2fYe80wVCJfVMljBFnKaUQrIWFcL
83GKOqJS4ecvjTSQvrMHxeI2Ncra0l8sqFxTMDEWstR0B+3us5nzUjr0MOu5//au
Hrh6a0LkZGwhpk7C4HfRTZemkq1SPnzRq25oOpOD1f8JrNRciz0z+3hI2G3h3Q5w
QECkFxW/+yhNO46tpcGP0vX4XQR+z8KdrgoFoO2qGi7NlIPuxcWMDEQqmIRdPju2
ceu5TcZKlfd/iU+/CY6n+PK0b5ncDPCK3UtH/8O33kTljy9d4jfa98U9Kavfbtm6
c4CpfazXfKTU9lIPohAXvPlNFx2iNcPaVNuRbvtbYPXrMOFQLygutV4+54wbC098
qpIXrRw6kHPhcKN3JmhEh6CK6NDTKApo35wXD1kW/mCALKvTcs+PQrGQbjN6AhqE
OMd+hKKA5LZkzbsF5SmQmMiB4ehqdaXk30v9C64OCl9QPCL0vxAbRhbkjXwVVHiE
IBMYGIe+E9OGAXyJaIKJaMKn48Ury7H3Ui+n+xW9KPdMBi2KpQSNAJ8RDM29jF5F
v5TDe0Z+eGSQ+uBPN0NLhOiISF+KcFo2bf5vdSmLr3N+WvaRxpJoEcKtyioAsZj0
W8S+F6Ag1Nob2VSxUJxe435K3h+llQoQjunZwa8RsWv0tU85Z8PWXe2m6h7pwW1B
/EcGA5U4keevHmbm8fpHLCRK0Y221KFM62Ek5ASWqDRjGkfOCC6jo8f6TOvyOc/8
BAr720rCJ+kyz8LSNLqSyeAzRWY/YU8ZXw0xuvPwiIuG5vl9Q6CWWGc43VK43UJE
WmKoV5kpx98h/SRKJHPYKd4i9nE8J2wZLUhxBvYsIAMzUBSfnN7x+UeQBYm6BXtl
95ygJ4vaPnkCQIUubdz4ASCbVWeqzJvUIfiebFRReeOeFRpr6SW85Xe17O+d/1Re
D5RwBOlGEr+6TlTVh2O+PWsZB5BYkTb319AYiKgoYA//NPyMeTPq6Rza6NhLIKMy
87sJwsn6HT460Fq/MA93q6O28mkHtwLt+1iB6nMvm50Ywwu6khwOY9GwuNF8Hm79
XfQFvvxHUw1PXvonG9Swc+zjzWhu8oaTj6b1LNTyg+Mq//IlL/dF5NucVu9F8jKo
svaCdDYFTsrkzgYtS3FlslvjZqHm3yj3vmEYrId4Kid8Rrgj3Hj3bZ/JVla7aHRn
H13C6AoXADUbt1DUr3oUMeqnVxADZAyrNYExOzhR6QhLs6+syrHM0oG96W4xXaY/
UWE1UnoN7c1BtTgbCAVadswKQ98Zj6HIb5uK6lgrXWCNgo+scnRkYwix4ULjPzrF
sIlPuPdcvEqQghlPU9ijDj5w56cvkftFHzVp1zoJHB/f8MdBYW7mwliF9Fvmv9iN
lV72vn3oy36yQ7op4V6hTGe66jQqIm+1ysHI4oEG4VWYRwNQkw6pDTuQsNGfYxyJ
2zRf8DgslYEQyJRePhXBqQ1zrMnPTJ9il6eYSBy4e+QVhBCUuC0b2z4zSYcBHHGn
lOlFOZkprsV3gHGcn/FK+YHNCSLsLyykNQi2zkL7TR3EDJo/4TN+c0EXNZDR0JW+
OiQxHowlUoNUFScRVi+q+TPAoZHk8HapdNMurQoT1wuZUjHcXwI9spLGoOO11RuX
xDbDz3ZhSodWGO7s9X88S3IobRCMXtnlft+GXJuJZyZZ/VytIKJrVhhkpjtLi64Z
/BN4KPmArLAgRH/FZ2vbRmiJkqJQiczpaO3aPM946iqGD6rBUaA4e5oggMYmswft
8PjupQdp9a9DmDn1U5MfgeRRGzHy9VTZvUDMBajnoRqzaAqgEOXdiP0YwLo6OhIL
PLY/zWYUEFdJoeg/Y/pX3ArXwwf7P4P3BMCi/0WJ5BokJzMz5ZeEF6t/rZqEVlee
DGEVncwDe4gJRe3c7r/3p2e53aC2H5ujy+IpCxorhnuS0sAacPmj/KZWAcbuz39y
EdUBWPzrjPut8NlHilJxwtZ/NT6GGXxdhZvsg17DE9c0MKeCIyr3G+1UPZOw0laj
pYWkRLVJ5I6Yswn+WlLRYqfQ1v/O1kcVcdy0W+sS4w5aAn+k0YI7KWNB6F9e3YEU
CUFnmL4dePJkyngXPut6VusS4y31BNvL7DEwPvhV+UmpiKYDrAuV1c1+hUy+BMzZ
L6Bp//aF2bZRBSbaGAGP0qjX952OPiAKb4xMWWD0Tvkj/C5Punva7Va+BcRd95by
FIlC5M1qUdTw/t19ZnNGuaof579DMPuyhAiopJLxfPDxFEYmYi/u/JKB5uzVoCeX
U5HQ8YrDxw1hW+SyGrGmuXea8/ezoIRjWLUrbkM5lI26LoU2p3DFEuh8BRUFIeW5
JgOzHpuoYEkbAGeRJMlJfcp3yvwOK5I/hZ7MAAVYaZF/RlNh88CF4YPDLsDT1W45
Rqyvyq+NoHwt5veoC6P/d8ClzvdJLdZ+Tj11M1q6QGfS9mw6mv4TFdsm7oIkxAsM
6nBzs7LcUyt+K64Tc9iUvirZFzs7QY4lq2smN9CTd6zIfxk7LqzdP6xSCuKaAJ07
hRSOmDgPy2H0YrHwE+khpMXhWGTGfN+ZowcVC4QczIXqHEkXTsGum9lv1Qy12f4w
ZdwoeJVsVP7GPrV2YzcAcSJRZtgpiqwWJsIN/dWm15jy5mkbBOJnI2DbcKLiWbdR
xefcQUhkSsewpiuCzGSKaR6oK55WeHal3ys4v1aSQ5FoEKFYXLtSAV8QqsvXFame
Jrru1OkDoPqOmxtrPuFsFo7muYXkF4mE2TtPhCMziPppHeerHV9mkyKgoMZoyz1d
IAen9pGxgr1N7m3mF+1WNJ77y/w0NtI+JMrHdxTuzCInccxx0IGv6165475DsD77
Umeq7uEVMgohBdWxCUvWiDUkxI3TSifpYgVPs1v23iWo78phybJFFcNoF18mbOC0
00iRxp4LrhTQ1AQhNRFrsPac7832LrZq+Iyog+3Gby8buMQiExHUHMxV+pmBO6y9
A0WXCmh0xvaZFLtQdwop16h2+6SebWP5ksQy2gwZKvNWQ2eZEWf4c/MM6YMq6dWt
q1x3LCVcXornvp9nWr6ogd70fl7QRzcf5JieIC3BBl72N0BwF/M/HTeOOXiushcI
a1nzn9Q7iZnCz+gGqzUlX0EN8ghvemQDw1lldSOHaP1sXA9eCv5qglokPomTCIS+
4T+QhtZVocyrjKE51WLCJ20rI+3xF//EsSbT1/9DfgDVLW94sSTzZGqbNh+dFPh+
9o8Spv/Lt9KXKdadPPTI1prL/05gJ/QhV67iiXNCr133eprtW2s4g+Bq0FqGBx9r
GxXBWRVzfZIUQilxUBjIxxd5Rrn6FUtCQdSCL39+g8xWeNo8rJZksedERB6FY7+d
YTpywA9pDhwiO1Q/6ChBsr22WVSTJBt79VJxdg/Eae2SZ/54cOBuVzGj+uHq+FYV
oXnJQtCtHNKqkAHUqB0EHInLG+jt6LHV0k8m3rgIeBIk7HIdr6tlwYbb5pS5LmS/
axQv0TmdNEXs1aqkaG61iTFbvdOdZPGFdM+OQfI23ksdnKiKezt0yom++m4QWFEg
m4ZAR64XXBsVF3SEnDcjd5OIFDj4CwbEtNiSKb3/rI76kQo6QQ+VRlOLXfuT3Iu6
rMva8a786Ow8GsKfZ51oLLf4oWR4XMz500xKY2Olb7pqKRm/yogD6NVFa7cWlFyS
LUbb1Kyrv1D5fDAOAV/ETtAJWBenYzCiPkQhqki42mL+5Am4WxrZKxosK1nNlhkS
zchxSDzVlTxx08g9aHHUK6IlrDsQ7khbOi8ASTxRyFC1RZXuv0bv4SbXOpj1TWLn
qvFqLrEy93H9hVYrNPC1Q+OtYTWRu7KUC3Vj4ZRUMZdoX7+HxoIm+R14KzpvTY0m
JUSEWhqIpi+UFmRT1kPsw8S+x5Olj1iXG4FyUKUBbPXijUki3IFkqzLcY8fZzt2o
aphwEEuSAD29mrCULO61pTzy3VAXfvfgItZNtPdpkKcFf2v59g3UP5dVVLVqmAUR
WjAjLscg+C3yiREJXcPms4K6DgJEkER9E/xyWouwl3bKP/ljmmZwoKPDmKURgI/7
L9oLKK3vZWsizXi5ZTuMs4NJUMY1IKN8NJDmbRmhA6GWCJEEwidveKdpcDnL/73a
pTZ4U2/S4avvpawG4g1IWDOOROoYk919EGCYq55sWINxxNt0Sr1bEktsPkkPn4nr
W6N6l2b/ZiUCE1CBlhyYLXDt/2UwsRWiNksZnikrMso8XHeqFRkqw6Ep7wpZAmJx
vV0yck/pcJTMitwCnXTdUaIMNKbLeEPigSo8JbOX8Fy6uaEREIU4ndbGaT6q5ELw
agiYgBgYXQ+7hsEfZJnaq/CEvWpa2c+n4y0i/54a0lXSvFDWda0i/XhiteR7bFDY
Ux+nzsajxWvpfW2upzw2TTOq7x4D4rLDUOPf0uQZ2lP3Fdtsvqx3XRgh2tBUbEs9
4myQ4EdnCinbz3TN5dtMTk0I/XhDsIMNZhxC+/U8djoBxdqP+/SI5mqnvmjbsok2
c0sdKmBx0ql6cz+0OcfxVRM1CgVJnJU+GQGQNF4oXkK694wxyn/Qm7TzTZPu/xG4
LUIpniNpoleQTk6wI1i5s+0Q1/Yf41MUZ2Kfzh5lGsT7q4iDxaIAs+G1aWsHzVM4
Wop2abWOuoChzC12Ib9+rtN0GTRMZvS1Z892K10oXW3IG7JJkvBc51YHCi2u38EM
lPlq1io0fk/S9qKMxlBD1AddZIob9B+d/0NczuqqVvhmzXWP8hb/cPSHstly1Tsz
d6Eh41Li1URkLCd2ANrnCYpk4sbgnb57o7kFrshWl3se70wrLjQllvgPyqdWvr7L
lJVwMc5KUF6qplgBZwJH3jbF8vlnWKG7L0Uv2FoptjKGOIJnSWjSGNR9Fg1+J3Zs
QQPyRgW3G1f+ckG7T09WhWMDrBMb3eZbbemu0Gv/malDEXL5tKy9ShAnafsFlPR7
tQLNCI/cMAP6YWMOV4aILq2fb7ZgfEwkt3q6O/KZJVanNc2TDIywh4euMA0+cyCJ
R8TLVQvrMRQEogjm48gfGC9MZ9jc6i8kVk4x0mErgkJRYfnih3CEDzCCj4MJl8Ub
Uqp9ASvEKombLYSToCRFYzyqagCx0qI4Fz8W7OazCYYeZ7uqMWgYHW6Dc/0C25Uv
WGv+pUpwqmRl8KOF0zDTFUJcmx5W/RlErOTDq+ckOvYu0si1cevrJ+hzBqcu4MMw
Q+ZDHzNqKKRdtW8lt4PpLOXEEFX7oIL/zMElKW4EV12LxMLqdq7hjlJxUOqjJS/A
erSyYEaRaRpEs19WbUoyRy1GkInqEwbT0rG/lqYlhkTnBi8VYa+/SmH1e5pOL56J
DQj+haNr4nJHHoGLNn4LpcmOgakcakClxohIopr9kQGAoi1U/Hh5bcQJ5m+NlDzW
XLBTbEDS6ajzGaHI2XONHMSUmDIieFx5pSFuNmOohAPyq4XF2Pv4UG2Manig53Uf
Te3hdsiQHFh/sK0owtYF6aL+MXvibZY2v+br9fLiyjMm9vnaIZhwoEaWpLaZ0yCv
6F9ey8tPavbQOt6Uz45zi1S4rVXx8BMcIVb6SPbms9r5c9zK1WtMPAZqLFI/rCaf
TZkDv64g9qUVznJj21gueMVtpSBKLIPADoWvzj2im7tVMl8Xilk1ETPbnc3FYhg4
T5HR2MaVRPPdihWqekxzGnon5nkxWCt3xR0DEySvSwVpnulegsaBMvgkYLT7Npse
y71wPn4XRGrJNkPML4N9Q1uiVtVaVKfn8++7Aq7AbTSsA7vXKilY06iN4SqFgblI
lpuHPP0OenVhL/sWIADUgMrEZfso5Z7t/o8SddpU8wVzPWMJ2u9RtsoiPJwytnws
izK0PjnzE6gfmT6agpujsLpdRozIq5IWWYd7+gjlj8WNLrBuaOlKsA2bxEWZS9T5
Cl+fI7JYvnU6gE2e4sj4aTpnK9oVPOt+7vFU4sUiruyPXUcjQWuckK2f8MWzxLmg
OrIXLtpPlH8GEEVzGyqOKa9pB+1agPbvWqY90PH2HnfZV61ICf3OyuGDLZmbxrRs
yGdNcBMQ1QrRgXTX45F9HSpnkmLuEMhVgyVJfGnfFfceLGnl7cJV+G0cWp09Nhmy
uxj+rO2qHzkpUsM1b0OGM3SmtIw5RCLBSNmZSFnfoNIEmduIhQuV0TAh+uBZ2Xjs
1Xylw3K7l4nMXMUJkFvQ1dv5m6DM+QcwOeu8RyV15JMz/EaJdy83TjnG+i3kxRr4
sJcDKawx9Bcpun88LqkGfxoodpejgaZkdDyGcpW9fyePz7bxf+B8JCgin+xSaEpO
rlduBaegQPeSl4/FZd5P7Z4s/+Zte89O6WYP66KaPnR23p2LVr/c2ej1VPdOcMih
OSD/tqNm9VDo3arOYzgS4Js/t7NSwFU6SECAz/J+cCiEEQjzb3wgoGXQf9CaYhGk
fiKYBiPRUrSsj0+gk4hbP2Dh5xeAfF8SSvg739pbKTyEincqiRd4LjiOdF5tXxy+
wxAqEhzvCnkqZUxFVdKANivqpmRHEVKxmUSVZxwVWrSf9VzGKhf/RiZQzPZ4JydX
/WvIFh+uN9nrBbENvZMwWNos+Ihgz1rnIeFqPSdWuK4bq9zZgIbYJ9Zfpelw2H6F
WdJ7oimvWAX0b1FOq1EIEBBqUECO0iXqcn+d8ej1N6+CYQZyVN5FrRDYeT1DT6aa
S4AND+ZCxvayvQY5UM4XBJVfTZfj4RseVPWM6b8/6ysMRcGwGPHc8B95fnbJNyP2
A2hZJou3447IqZCypWqP8eYFXFh0XRR2DQm9aI+1PRPde+8JhgkVArE+SFPrXAcY
Ct7Co0dDKdJQ6gZeP9VfiL6BtR/S5FRbm8QkPYaRLVOYvUXKLQDCCs/ZsEeR8Kn1
H7DaXPA1C6C9bz7/C1PO04DYCO3nnZI6VqWSUnWAtTyqF3YtB8b/Owmrm740FF6L
B+UmzRltHQAyxxw0l6usNRZtW6QmmHyGrQRCnRvi04036Q4J0MmzGB3r+Ry1X9UJ
uuhTBk8GwFjeSfrlAaOW7Yu3jl4ABQuMqR+8XjGGlpozonbo8PUYY8/iy/pXUC6T
IL3ge181NcbN1+U4TdLZv1L8G3bAL3GalOL00IqhCc/yo+b4dXOk+GAOkLkci5hc
e2zphKqfpvrzq795ob/Lw0deFWrTmb58mfOc0tV32YyEgYpgUheUFP0tpl+xHwHP
KAOSPJEnutXIL1coFit7sa9rGXK8DCczDm/dL1glhBoKegH7Eirscg8jGQbKVhmx
o57SWOyeI6ZDXTm/VReBPHb1A8aPAMpREc8LVfCo/kGtXqZ4QQF/lS1cBsN7l3r4
6++kG8zyDoyxwMHryIA0XKV1qLGcNwXW3qLV7HV5catTLiNLe3Um8+n0yn9h6Ii2
AVH//YVdA3RwDsd2vEzE1DXLrCLjMkUhsnaxY1W/U2khCR0+Pxw196/7XuTAwmcX
fcU7CwWQduJ5WFhzSM/swNLDCyYY1u4CrG04LPi3VQj9SN6rGp5jN9aGDB9j1RgU
nGlj0QVxU0f/ZsCIxTYl3Jzu3y740zYoKwMjnLtDr0M9VYpFqFKcg05qJeWkz4ox
S6qZvI7ycZx+QNrmjqbTRueSM7TdPX711bhozGTzxD/GkywcVM1zH+x9OIntT0pT
4gJgo3J/80K6XnRNeUXKepVf1vTOsNZqLh9HlKSq3i8MnKvd4ajzoupSPeMSN3X2
MPaKlNEpdmR+WWhpbw5OUxMRO96jAdej5OUUwHxmwr9DZvDvSEdOER9uyuVRgPrd
4Ru5/0AgCuKSD2hJqFH4uLt4eMkr6i71VzC7o7c2BTejTai/yMpBtZkf3inRLWWE
KCFAKkUXhBA+YxkgFfbaG1vnLA/TUb8QfX+uqZDVw9nYa0DKyicWywDJ37Eey9yL
up7s/mMiu2CM74MtLf/IwZn7No85ek3+UFRaKSiNZ3skC+heP1LPUKyL1Pv3mRtZ
G/1Nag/jXZuGRFZBzInnPhmz1yn0qoBkSQuV+AklMZjC4peOfHp8c0rECS/ISVtg
bdFcMUwG87yfl/tSblUa4T61N17QZDpRQ/lv41Szu5LNKX3Jejy2Njgbb8LyIXGZ
gzKdNOd/sxWoI7USZS7V/7PIVgg/ig030VlVAD30vT5r0QBNTDWTGombK/ebzsWx
zf+M3Kl8qGJA75RlcITFIMey3jF96qDG0mcHs5yEBx+lHeHYgaFMgj5J3/iXVEPD
HKPnW4WGuAlBYtwk3rYVq5vhGUgSV0Yby8NKeaumHbQLbj3FrePHnvlREiHgTqG4
Zhh+uSAr91C2/862N3SAIAx9Ah6nrHi6681qzwzXldPj5g6juOrduiD/01aQRmbA
7uyLb1YheLbthet4SmcfTSy6H/IhnCazo9EDAY5/gwKlKYs54Yqh+tlwu1Qk6Wb3
+wNE5G8PYH5IRebrgNP8u6ypwnucB9Unou2F9iqU+gI9zrRW+47zLaH9XbtnFsaz
fPf7ceL/XTGLQVdHMw/fpMi7EiywJW029t8/9IdaP1weJT8ilX9kVzpIzUR2UzoS
Uw0Qy938U2ZQzbHS3T74wk8ELgEOzB9BboLSRDoyERjpCsznLRVsiiFlc0oSGs5h
101GNKE1ZfHgUlbhtfhG5kc3kFMYsONCb2wTe24GodgRuiEbQ1bj94ZyfLTnuqCP
7f9+xncbkkJD30/4mv3rw2QjAAeZxm1lDcvYfdDvVk1VvP28zDjUUOR1BUCr6zsU
+mUoWlXhM+QUGKqFOiKeZQjebG/+XCpvcSCWjYcKuZUtxcA4aaWW8u3mGKyq75UR
cbEDMEXTO/kkcEIANW99IEt685PGMLsnRBuX+TLL4DtVJW2c8OEqs8r6/RQBmL2c
XpU/biVkO8lIEuqt6hRorcDLySUvEPD7PSs8aJSBvN/0m3GrKwp+3C7cjmse0pkc
jodtkV1Q15VWqzuYiIFrFojXh8xYKJmhpVmCU61JShZ//ULmgbRlyX/ESWAm8fMp
sv10FjfTCDkqEI2Mi4r0DDRFWfw8ADjX45meKN1yoLe2hB1RnuQdCXzWsfbQvYCM
f1jq+utrUJkegaH0YMr9fQ==
`pragma protect end_protected
