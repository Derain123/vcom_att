`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="galaxsim"
`pragma protect encrypt_agent_info="https://www.x-epic.com"
`pragma protect key_keyowner="x-epic"
`pragma protect key_keyname="rsa-key1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
ERDV+p2OhhDt0abwYVgY4pb0HfcyndhZquV8+XMtxlEla9WAiWq+pZDJzYzMcnLo
bSHSWo+JO4wiS8NdWHcGr506Mixc3wb49PqFGzOAHW/f6seOJLrIa7bYFBEYnKdN
YZ8MsX8I1Ua1/dJJlQ+OhUTRMIgdt87yx6fxDyPeHJEJr88cnrd6jfyqN/vGEaCh
Hj+HF1fYRU3a61ahYoW9Kw8wjvAbUmLceEOw1nbt7mwC3XEjnTDnL2aqLp8QwmOn
9aYdMYMsliIFBG6gu94RnryptEFauiB/+1zmrxTO5hzjaA8yhD12hrndnllCfVJK
6XyTZomhglGwOyT4twbmCw==
`pragma protect key_keyowner="Xilinx"
`pragma protect key_keyname="xilinxt_2019_02"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
nit/ChbYK0xGIKh4Mr9hhosd2Vo5bVvdonykDQCr2Q5RaIZj4qfxSDUBGukbPWkJ
MNzjRKm/uUPf24G3XA0S0IRrG2mvUjYF4Rn5RuD0yli4IETWbCsPhrMQBf4Abrxq
y7J3ShMzfskN9Fotn78lpi1VTUVVH3QUqRyfP9GPWgqSP/IaFXZyCrQ1RBHh4H4G
6iwzHVOHXyqhIlduZYxRDEcn+xGnH2pok3kVNDxHWClpa1SYCWbboa8h3EOawAiP
pii/EGCYQk0hsIDdo/p8Q+KObrYGaECxXjzq1LUiRyIzoD+IpFKlR0nxdbDZObLc
CJxn5W8+i6zAEGdMrr5oRQ==
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`pragma protect key_block
SppjqKFsfesvf9kDwrUeWvUaIMG9X89BSaztF6MYm+PcJrTKd+ZgzjiFuZBtoAjo
nWxJNmDB22AR+QsaS/+mRaqYHavT7iGAutdgHBSDfOkqpgjEOEJxh1oDbPN4987Q
0B96qe/cT1LdH83dnu2qlAAyJd9zmY1soeJhUaio+iE=
`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
S7Fl3ZuqpoN0c8Kuk0jaXK3yUD4Lpav7196gBXK//vZZePeXnEWdb/6lCj00Zl+V
qmJnFLNSgRyi2cGvK/8vo1XK1qssv3/zexLsf169qAOHQRyqC0n+5k9bcxaI3sRr
5AcdVoCV0sxzrPPv2mUMD+/Qw2ESkSJw5NJz/h32pvTkApW0yyXVTDgUPBxGUUlQ
AYcfWVoS1ZdYW9hmqqEoFtrXvfeidK2M1OYyn4WEWY4rWzl3tTDlEWiDs8/0qY5R
Fo3WlLjV0N2Dj58u5f8d+OgcZjbKom3vwLIPTD4cuWbl80B4hTB5NRYCR0DBV4hB
XaMhLzgD7DeB6DkWPdPA7A==
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP15_1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
tPbwZA8eWk3BGeKttdOqo6xbYaBO1uipFWsvx6CHgJmgjrkUzOEFJWpZXI8MBq8Y
Kiurrj3kcjGWoAU09D1dlEmN0dYwinAmJtqDeuI/3b43vykL92wKsgy+b3HDIsSl
NOqutq3rI8ug42icYOPAfy6XvWNc5JAeLRNo7UDA//2/erslTwTQ72gdvrQKyW5U
bkg5mU28FFPcE1F7vKy1q3WO/e/9fGuyvAmOSY/2hN39qShCeGZmkUY8RjjbtYWq
pRGSgqeV10NLQFtpxQZE+lihZOrrwz89cdIiYSlethvVPF40vuxD7QcIPMtVJZYP
R6t0d2Qic1/3miHTTJPwTQ==

`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 4944)
`pragma protect data_block
VP+WYyxh3WZA+TRJEmQuxIpgzFlomyYxnT1FKU9QIqMvIFKZQ3av+32t5sfJoxTn
nsf4yDjhuGEUzc8ZvMLiKscCvqAgVE4pVzLuBuGJfM4KzZQhprARrhXFT3qdpmQz
9fYj7Rqwlo+mLtAvsRBRIM8U9dyoj9ZtKs8SPlTgVY9jb5gqTqq8P/rOmIaa8gQr
fK76kdZj3yHbcPmVW69IUck9SmGb/yQH/K7hy6bJ6FEdBYbI0HuQ+GSvYWp7Iw+7
kykyhe26go2f3gefPilTOwjfKjLcsUqpnfCESQLfKTTlKHnrgPI8/Op43ZckN3s/
tzBZEri8P+2AeXVtpbfP8vnU5RO2DkCMdrLYjMKuGjiAoqG08r+ZBiqc3q2O1OVc
6SUgOYu1iBEKjImTRJ/n0ovATFD340uYo16Ni3qbdv68aLbf88f6gx+WBl4NGR0p
80Owd0Ry/4XjdMzEwSPeRNUDFZO/enWBGNBlNedj/UWPcE1PPp2CPzDIRj4LoHtn
QeEjgaH5Y7VgRHLvsbnUqpAxfuD6Oo97ffCrPzGlW2EO7ry7SyiItzma9BOXsrBZ
stmzYLwEj9MStSrKdLP4yXfUS3a30zOdjuiyqqvkBbkrSDoRbsGttj+ju8biTg9M
hO9lIVs4lGc14wApjD6zkHBEwu+jQVOG+RYrMK5xXCWRJ4xqGbaqXBwxcgJ3FP2q
Vau2QhxrkpbH1tTTyxcVy6Z1kg4l7W4jHnVxYX6SBTcgcMYfzHeaRkp8Qo3UKK6r
w8eY0bTH9+qKCrjsObm+IfIZefDoPNV/hRl8H8jA6NEErTawKiIYHQP6Kh5Xf/p2
D4mU+MZrA0rv7jZDS88nC1TVC6q6VezIhOqXkDcW4WTRD09vL432PB7u+aGHefNv
kmJYsjNHMBEkpIj3vITcWqPC5NvXY0E+G+DYduCEndhxTeI0uHMMw49WaCvlsnux
bhtH0vMUxYVO88y1CUXz1EchBSY223J4AozLeOsy/UU+DwejfY3NLBoX0R3WffGc
aFbFi7anH2nU+JPk5HqWlvNuqXa/krEBddgamYT/Tf5lZZJ4+wu4i6OUzkbkJRi3
Da2o+mdVo3UNxihytqAA2wrxh/LlIuv3Tq+dpUlRO8PClKMlF/qvKTlTH02S8tBw
7+/WoAP5hvb5a77WoJflHGxRqCEI3f5LShfBu7qEP5FQ0QfqdO6Q3CJodEaDvf+H
32SQqM2k3JqqqR0uMNnx3d+z69WLNbz2HSY2+01++Il8St5Ev6rX/nDJmcI7uvFv
juYDPJx0LfeYXgMFK+392Z6TAMIHAhbeOEAtCwZ1pjG8VP+z/9sWf4JYAPXClsVd
gw0Oi8IazetcH+Hw3S2CRfhRmx+5dZysHa0wCH55OZ1xr09EEhh2QPvGrRz4Kpic
Xg3XXFmtyj5WmiavoB9hxYmM1tDACLxeJh3SWsYxZqyrjgKFC6YAJGxcS1SbeJ6/
HqlRsJib5lmaZxLvPK2LbHRCyM3gChewLK5rdprKmk1SD7mR5SQM9JrBPM+zjMlI
4FUK+Kuo9qq7ZTYi+r4dNCD6YEgycDpKfrb2RU0oqJGnL6CeoqrV4FEcAfbXcbht
kPr5krGCe+DvGaqqNb/1D8e4loSkcGhfWHs0yP2F5874Roaab39mVUOYqz33WcYM
gZdEOwmr3Qvm4uObu4rPIVa3BUozJyDsjStqmQlCpHzMeUL7tfm81WO0nIhu+WDQ
STgB+yuOuE6Jt1WyH4YydIXjgO9FiEMwfYr7ZFY5koaOzjutgw/l0/ZrXmIH0xQn
8AF3YAV8u7qsEtgRB+tWrDV+ZZG0utW3oYvJKIdHukMAUS6k8/BMIR9eTeJhvWnP
ET5yDLlqo/B+YdSCNd6nHxjvIoejko4vFGcJTDoe1nj2zizmetSm/zClJf9QwrG3
t17T+qWDFRssso8v8+rJxJqt5AaHJGDS2ziw4AygaMFky6ttDgaplZtdtXCq03P5
RSYPRHsLxKBDP1IxMfCBn/2uhQ1hge6p4N5dTYIYvFJoVaPgSDqrUuR7hcga/kTx
LULg0ggR1PUd5i9emlWFpd3c6XmmZ6YgMvFiwYMVoL4i5wni60HFTkTz7p6IyLC1
tGhxHHSrYFWyuv0ZmzlWE05lKWY+OgkhxVryLUrsd03jDOTzVh4WIhBza091rcD4
kykNSxBsTpMnLzGxQFSqbtwY4usF+AkoFiUQiAMZgJTAFs4kcpWrstF31mi/ellV
no5caB4SABilJCINCME49XHuSLo/KkO47L25EHtPYcMCN0U0c4yYF5X7HgKs9vzN
Fg8PFyik9J4/WVnJf2VMel77r02AG0sGm6X8uVhlptICbAMvG1WHS9vcnjCCba6v
dqRXnJylBUL85//QJJHHqjpzdPserkPeTaDg0v8Mr4IEp77Cfv7X57IryQzpEcbK
+VHdGuNoxhXCRTNGjAzYL7jrrqwv/o9DzQk4k6LbLTmC9LqV7dYhzge5Ebgso5X3
H4O3QNTcF07qnkqoJeZi5mMmoH83SuoTecQoI2tgdSZe9gkHAlc99qe2kL2QAcpx
6GWx0Rh8c7dlEbyoIHdTwu8PVvAnGvOBZ8rRAEtoOhgw1KC3EPrymdFFe/CrV4yu
7GbNjJ0HnNyg++puP1jPw2cw7ja+6QTlq0l5Kk9eUlJy1+/FLuVBxvHPK41B9SSS
RTBbUd3FqTTHRpX0wkiyC8ZXvlkQ3nymZV8v5HpDOOEdmm5DNAQ274dE4AzoJaeB
dC2S/LzbdAjDWxmO26I2wrlBQIp4Wi14U92hqx12ichlQCWKU1vyKX5VTvCpp5OV
d9ZvO1Bwg/pOBxjvZNZkObC1IBEcwgyYceCdggFPpwlOX8m8SQahmJNNzpiZPu0Y
E+jQNzm0JuKScWNTDFXus4EaWZoP23/PKyBJ8mxpFGVLnqJzqdGp0DUify1Fugiy
yghYHr8mALiPqrA9/RJzkpr7GLw23eqDzrKLc/FljN1uzpBGM7aRziJW5TVdDTZn
7D7RDdBB9sjCYTN7rVvYQNmF/GwY9LskORU4F40bQMvrb/hdHyoQwYgjf7iPRsXB
SSyduWRYg/HQIEbQD9YkEgssuBYf2/5UQGsmDk8x6dMfks3R3lb+xMnz2ekzK5NC
v533r2epCvSEHcSxzSxU7/xs+RC2KeMQQdQxCvPtKQZamyH7G0gAFCgMpDdMHR5B
0KlaSq8PqeUKrY+Q+WXnUAWZF78bt73TnirlSsWrc+LZwTQCm067WP9bGkFrxD7h
1Eb778wNu080ZUOWL8CDKRqNkKG6+415ez5dn8oabTvI09v6mqjNbJOLSktGmABw
40A+RK1K7GnxMSErtUl7IUTRBnQNWMHFN6ogQAE51XSF5MawbPv4Ro3A6VDU5Zal
KYj03C7TY1IMp9WFXSNe0SRB+ga2e/itdzl0Tw7FGxmJ5ZjcYwuKRPVH1DMFQmEf
LxI5ZdV7dT5NqmH6JTWWTBc/4skV7LMbOhL2n9HjvZFceAtJSLT0SbHq+APSi0Ei
lY+E+yqh8001PN5L+Nh/Ciws9RZEvM3VIO2Dwi6lyHKYu66GM4bFWn9CqA0+BjVf
mgAU8ddeC82EasiDDTKB6IGFs9+AUsUFkBtxfQbyAhCB2TxA2hPJOrM6iFNuO575
wMHs0Lwm+nKx5BwBFW4yty1KbS7Q5NZDGwGwbRcUmm3zczLb2u5/Qz360Y9+a7OQ
CSJxpAyoSs83feiTv0iotyTiR3UsobtnFvV5DEf+9IA13TBp7yDXyt71Xg/IEZCH
y7DDwtm94p262caeZJWWSdA4Jf0rLkmSukLHaRdoOjMuQMmpoOUebWHWoNQgNjex
aqIvcV65BkRAEo+Dy0WHzdM4rsdYt4Mjq7JBmrT5j6oc2ehnjU6HBM2yf2BBstXr
+MB+RGr3H660kjyutNZOwjOJu0jH+pGNh/bNAE7x2Mk28n0PCQqDFRqT49OXIqGu
1Cc6wVm2s5B/0EkgZQmEl+galigP+IV0iwMV43o3oMpSqQwxkaqIOXfO4+taccOn
9vZTwn8iyE7qdrbVq7OCT5oWnaS0Y499kyxmGVuEGiKImGpzGb1acBDkg/XuhWIn
GydEbYt1xFGGfiMOKLZ/v0pZtrtucjfcG4pC2CT/FJ+ERaajXOHz9aWr+PZ6kdOU
lCJ12bb5s4aQGaQj2xoGkqvjX6kT3tNxhb/PvX8EhS2lpJb16xCeyYfurV8+Mwpr
olvu30RB0GxrbVPfHafcpl6k6g3oP8uNr1PQY6yYQKVd8AjEivCfkgKrsxIQX1ri
dprlC40aIa9hU2NctDeYmTHHCodnVDtmAgerhC5fRm0nzu+FuDYw3S96hvGw041G
4V0pV2WYzERInW3zibepWVXgezGEY+E2M+sUtAOX1UPPx56SleuYtkhAI766DPkY
+GgvIhLtc2833qd1VSrmSmBZz28BMX4k2nNlmKvwsYWrqVRv9QCG110W9fwuCotb
Woe5NeA8Unfl45z+RLTgEuRHgiPomgxN5BDsARq1pFMKrPcx/FnWrjXa4E6L40JF
2kWxG9UITDg/iKE4ZGhCA2z5TI40dE+qqjyrQ++EIoMwl2r7EJKyBcaCEfdyQ/2f
S1vC3BohUTaTFVY3AN9RA9Pqx8pXScCQUoePBwGuD3SCgO6Ucc7yhdkZhfykOR9P
lXG3m5qIyWU+i+vPIlTnKEpUR+iOi73YpDYQ3IhR/Ur/7QTzG0LGI7Uf6vkBW2Nc
SNIajjs7I22G6sroz7edtXZWL3Xba7bEQjJKRroeNDS2d6eJy76jX/lHXkTAbAUo
RPBnkOwHtKrwC3z4eQmWXdLrDLXNSQshzgSUmy/i1VYgA8k0R75ljHP+ZhgNyvwj
uHMczmgkogx3dd03qOlxzYxChX1sg2Nf9fEU53O8yjFffNikuAnPlO0+5BduJb8m
4phCDcOOACB/t98U4GeeLxvizfwMqA9kFWWllEbWQAPZEuJU/Wzr8ft3zotRku6k
mCz+qufv7um1RlLrHM4ywjYuQvDKEHLDs7KexEyfiM4mec5C8f5nOAVCh0x0fRrr
G2pWdBUoVxyIYkiCJLfc204p/sKhp9TEsKXWZA3OAoLbLvfV9oHpfbOhHTO+Hght
yS0jpjFpCJqQ498KWtWbVSzEptgmewxwP7xLHoGPO12YVH67VYKHuIKmaYz8OaEb
d/Hq5B2jIvZDO6sUuh4oIqCCRv39g6U+jJ6NSVDgt4QiEiF8YonxpA9DFJLwSzLD
xkQxWPmvUlzc/OAYwfKfonr3j1s0R3fUuAKGsgvR3wSTOEuaN1tBcPIA+q6s3ieH
bYuzkTYFKMLHRTcg5iE+q/dL4YnwteJ3P+ASTNI6v7gL7LO7tsde2Xp9/Sl0I0VS
Lo4NfpfrzFOSSRYzZlUKDeH3C98rYftbfL1Z+8g6Fis2c5gY5q4KkYDvrPTSbv8D
wUBkF4Ec3DsFYhqWdiOwDC2vw1smDbIyLrP/QyLuJGGedbITsoDvF55/FVwlOIvw
3qSt4hp226Owk+6dugyH23J2iT9WkwDqk4D41kZ9Szxc2Ob2ICWaSz+w4VM2Bwb3
OWG0RpD7MMHw67Gl3+75hhAQJcPS8uGEvAiuTdWwFOH6iwjTl1lEcOhDWJJRcyEU
SlrX9rvKqRYzLs1neghJupFJLT6vTPR9MTr2iX1wiOwH/x7Zl+xKiAj8DgKOksdC
ddE7p06uDkCBoC9KbtpNGtf5kP+0pMBACs8B/dcuWgvwETAf4RKlSHH8NTqLKQep
Pj6MG0C+WW1AzN+uGG+RASaf8psB/E1jOWuKJbG5ACSZ2dnhVeJsOXLV4tYSNJu9
ueJ5lAUQbPN3QoNrN3PYxKo1++xxtzt0NnUn60dpiLZW59ZhGkgzV/A+lRJUbZ0V
iShVuUMDatGaLhWIswyL8yRyVcn7NoolEysQ3W0I0PB4k4KOZNfwV39ftlxK8wU7
EI9+qZOC8+wa3zxK/op9o1+ZKRjDfGKRIbDcj81pdxQx2RyPFto0uzba+Z8Mqe7U
178wSDnCpeUg8LjmYb5ZcYnr81Y5pMer/Q3Yxu0iYyF27778VxNneMZvAxhiqC57
/j4FF36yLm+Sdphq5OodZVoYoBI6x0OTJ+maWQAlc9ICIWEBc1UlnmtolpqyVhHV
NBHno36AbkWLd8mUDWPL51YBcnqjPMJasBTGwBmOZ6e0vdaZWxPS7+MKImFWajaP
0cWySFwx7IE5kMXPgMg+qUMEaxLEm6TCsTLrqbWcMEEcwYrItTWdC19N56vtMlwZ
+D4+MGD4j+49jSob8Ij+naMXKcP5CKCUU7ZRIoC7fbXxV44oB4U1OxxOjfhZbOgu
cW+KvKntHxsiJ0ICwcrdoV/48GC3QyvADCnQTJTeFn6BXo/+vEsYiVDwyuwyUMtC
lSUwB3Q5sPyZG8Z1VQpEZp6X4BdPMqY9Ba2hJVQjn7pgy7zVuMF3cLhc498yFJ7G
KonE/AaFIkh54wCnLPwc4qdkhPyD50K6pI5TkfPOEBzCSQK4O4NlCOH3AulYySZY
cMpgW/54UCIXzERb9uxEMEK7l3B1ZO1mk2TkciV7nQKL0UxbPCkUZhAboh09BSHT
`pragma protect end_protected
