`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="galaxsim"
`pragma protect encrypt_agent_info="https://www.x-epic.com"
`pragma protect key_keyowner="x-epic"
`pragma protect key_keyname="rsa-key1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
JRTaQ36Ve5KkJ9yXagQHYOwavqOzVCB/bQDttlm+riNZoppv1SdkXSkGfdWvlqTu
GFddvhUm4GXAveWPQ+ACTtjaFWKBtCgvog6M8QqRKJISQNtUHk6TgZfx40CgRsuY
caXoa8m3u96L95arsI2JC89CO46CfgNfkBpcb8tWHWisRzjklo5ERTl+9GijsJQH
2Dakn3bo2bqEuedKkDZ50eY2gGbh2WxQpHI+KoLFHYpbumD8OQfDKqSosHsyLEOl
oYxQp2Ol9o/tALyvDbUYkCBWZV7nid69/3a92bPS1TmXgOpELE7aMuC+Ir7nTz0H
lXeZ1RU7wambGhf3Nw2DMQ==
`pragma protect key_keyowner="Xilinx"
`pragma protect key_keyname="xilinxt_2019_02"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
RBcin+GpOoW8cVXT3C51s0fMle2pupA9iPENagpldkXxmZUGADhAeIuMKNfQS9Zu
hNaMN1/7khLLTy0wdyvmo3iM4pxfAMpT7j0AcKoEGHZSU1WmEGNeq/smj155rUyW
SAkxcdasbEDFkJqoMcznsrsE5h2rZj2/6UZnYVzlhSX3asRj+mV/z714omzy5Jxn
0KGUikKAs+CVVqw+zJeFb6UCgE09W8MfT7o/rSnKDPixJKK3jPVnKL75jnxGwhMv
tBMRcYyj8IE9tz/R64PvCzBACH4I+KRMG6OeLvDLRc7JtA0Q49H+Q4hHm/ua0LhM
r5onKID+sJKl1dVShNTj7w==
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`pragma protect key_block
qnBL82IzpjbMAkn/fC0N8ulaREwqp5DGq8tXigkvCJk2/rVd+KZrIsdnuEYQ24k5
NReSUc5pD0hX7eKBXNDnTwBIpNG+en3N9fX8au6xUEvhCreY8WCA5rdRNw3Kqa4n
dMmwryBkj5ejU3A8rpgA3D3MlF1c+kOXnmlqr2ELI8g=
`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
T6Ah7Hv1W2njl7+qJsLkeVCV1f2lImwcwI2PUYaEI5D21MsQF744U8VF9lQpEVLE
XE1oYzFnjOFjd9W3XzEpYIyehg/6xk+NbWJoqlZH5NvIpILOjBGmgUfmYtyW/Xy4
4Koy03jiIFECx8KEQ9PG4aIslnW1vihneGer5M9n50KEx93QaJc1/6BggKFF8z2x
+hXgL6MVuwrZNWS8QQiscq4v00pd2M+YTEAo8O+tP7YSKy8res/6xkg2cmdNVHoC
Go1gMVbJYM8XVyy3Kv1e3skg76J4yh/Zibplc29vG571yTFJO/Qb/YzDHQIB2nNU
E9oECfiV5I4DB0RlEuFIwA==
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP15_1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
oMbPqBm1uoP/qthQhxMfWxH0ey1CZxg6lKwdsPSqrY9EXjJOhr0Gva8T7ZpR9PjM
fcMgqzCcb911YNZpw4F7R4FuHPPKKgl0IGJGGDKCnvOuJqfAju7Fz6WUCUgvEGS3
8pWE9381/MLX/MaKeahVhBVA8T9ziUY5gBs9HQ12nMKcm1xiuKK1B6VecotvpnnI
IuDP3mpEb47jXZKvAK1v4YsV5C58zUVPOOLuEKz8S9RNOtuzFKZcg9orVSOeb7ud
50LRhggzIU/ioe6wqhx+MZCvghEQjKNotznhs/gxjI+C8z1uAUjCAwggM/AlDWYl
8HvGWXP9XQpkpPmTdVcnhg==

`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 3456)
`pragma protect data_block
NwXiMjDHcObBpdscnrIuj9aV9ckoI4JAODZGocH0CuctKhtjx1O//IwV3a0ocp2G
YbJGjKAJ3TjcuzwgJfXXvFAaCGqs9szZuVih/MeryCiYuOSkOGFrgg8LWeZ5/LMY
sNxw5kXz1OMzHHDwiRJPnYBjmMOTICO86y7rGweqwCCH5pUzfaRSE8SN5K7QKkJi
GL4L5dveYRqM/2xFBv6ulTN7BRVfpjk+kA7tGybKr8U+Lv414swIS9ck+83ggcma
2Vjn+ytAPH5I9sjkGWSHpCa4Y72qKOtBGwW74nIsdH0N3B707BQfoi6I1W763WXR
VR0mJNfAPCeWMDOZnDWv/B50cjvjZWGIX4E6lLI70FCdtgLItAvcC00yF87qxGiu
Agn1kwf94gVVFI8tiXwiLuq2s2bO1PWAoZ4Wtp0wJWx1gHOhteMF/Fznz5T+mMal
8roZ7pc28cj0rsxgsmHvzSat20QPc8WN+eAljN51do17cZ+COwNW2asRHbXAPrwS
uP/KY3MXV1F7fa4BKFeQTifQOPr6mLL1DnRY+n8+vbpFjq0LNW6lFPo/57yrgdcs
LFOJ38iR5KQxlFDXYOS79YaPFfCMdUhPTg+SBb33YhHaZeFbhY6+Vw+zquFFsqc/
tBEEL5dhFUoHAQK58heK+IFoqj8NxZ2xscgHrxMfqsG5/23Lo8PTiogy8n2fciCA
DVKkyE0XkthL/uyq1HHDipZe6hXEfKCmacWSWE14vvhiSwhlh9jSQ+cmo/yji9OD
wpdgLEiUeEx4HwspDdPL05sewMMiB8iYw8kHNL1LE7OhR7MU/ZsV03REbr69v6V2
O0krrHIXfci6KIgHzk+2IpyaHP8NAMVn3X4ITs5hJLgS2SiRGkkV5wTGxibh8VKP
37NqTQguEh6bVPKn/UyDLBnmrtjwOgut6F2q3w8GwRfvFM14WOC3ZMdYQz/Jafmc
zUit5Bf870EwKP8Dv0q3SbM66CY5nRBWd3+bfndrxx29bvYAO7S76ys7w5ExizgF
8me2cwC4NGL18XVEbHVMr4rSHXViCJJU86YO0+X7RbO3PGbUW6yERM8h6jDzJRNp
Jt3qVsq+a7o8q0zUpLs8BAxJGKA7JvEjKxY2mRHqNCEs2ki6cVtDY+StKba/U9YT
xS0n5++ok2StBzmSz5DFRJK8oBeQO72tGvOj34vnGdTdpxRyqGF6907b6+HzwF5C
I0ULNNL3N2ZUGuzjBp/Up2qq8CxWjOjc+AOalAPZFtZcsAISMzfKsuCgEtE2FTWr
RKKfryNGmTVjYj8eeMpcoehPYfTVjnpBmkEgdWcZZwThbZCgIt9oPGqOC2JQtTDR
KFOQkaKz6FWjYbDYPn1JDUt2bNFrcYwWYjAjjDuHh4Gxk23aX/QBxR3W+iPgvevL
mzeQvhbtWhmyQZCxtwJjxcOPGuzB9NSLaZlV4UMqZxHHpWPYlLZ5olfUMzN3sHod
GlJZtynXnRJZaGLjXU4Nq8jAiFUgNJzYk1wu+2wbjT0ZIkVegF+nu/B13oOarXMO
qiFtQnEDqmvBVuiTLCLeGP0hAfF9Ii9D3fUwko1h4X67ReuUyvrzXWEbF/PGVxG5
M5OLdSbH58T81n1ZL6lrmvv1KFWXZfpSGetQiM1ZXkDTGgVJnelSmDJmiiWCYz/V
NTxIcYxTbDxXwOXAqZCVg3hSm3N4oqs6ZYcNL8A5B0p9GBeVYOlwZUhaeGnxYfep
UtMddadODeWJe8nCSBQQQlBJZpgwrw6JuiqSD5s85rmSMHbsDoeX0wsoR+HVA13n
CzdA6yikcWQ/YHusJpJDwZBs5fs15GLhrUs5CtFteOseEsKUVlq2vUiPWcfT7mzl
ukZ0WTjLOxbOkEn0/DlOGNyRxqZ+gEGQqVEOXUSvJ5PKgb3BXaPFxTsfpkAD1WE1
4C2qqilg35dBayNJV1d3KVdASMkfZkKU7EQoIfrANmksJ7oZufXCxpJmsYlan0q0
UBtl8mwsRW4Jo+tLBD/qFxuZe9g4vma44qkdAoUt4mfZ5uwqoMGC6v6bWbZav5hc
9aujrukkFe7WGD+zQGqb/Rqrz+jNRD2rPkqoeZ2jkalw1ibziGaPSd5wtslgG5pK
ISu5geFIVREM5hE6OvZ9CC0iKXezPKAR0LMq+cvpj4kcKcR1hHMMdktJkxo/e+6g
NZgUoEogVfK6dyC7G73oeGlMuTiX9/S6Ao+cadMPT/yPcxRvzY9vU0nfx1hXXPrO
00AVrk7yjT1k9iDtaG0fEA6m6KnYhVKEX9CqP3BMup/I9bQZMNGcI6xAu9to2WdL
N/sSioWU0qH4z7B6VmTdyWbxM0zRa3DsTqv/7ukGfjfhHnW087HyaQQcnvsUkYVQ
8tXXpTDqNwiK5xWz6ta6gXyUMUoOhBc8HWT7l9ieza97HjLKF6D8EpBj/t29pbkL
kli/xL9ThzA5syEdASJEooMbmk6hPix0NXeXCmLKafuaA4TmOYCZopskaabzSUr2
mYrZ12ElpDkiGWd2qGjLVdal8kLDVugcK1o5w2xLj7N5c1P4ShXX4NXP/sX1q7NT
tktXC2zwviwcInzQvvpL2Z+P3/kqTiK/2CQtUH5Tk3bUPPbAHpyzspLOSKm58UhB
b56C3z6nRC6QI43vB0BIh8My7NTW+xPlxUsVrv5zM28BgSpZ2QfM/9QWRLRHL2qv
TLGw0duw6UcnoJJhJ0/Y8UYSb+EKTbxopMldT3WJEmL3PPO/GrllqmxXr1qAv9lo
3WFlpYUqzuM8h81ng34tPexHQDem9XcECEjvmJx2Y1CQujSrth6XQ/ioQCP9cq+k
0J7LDFV0xqCsh93fAZBUG9Y9GS/k5jfS884LVF3ABuKjjYhzWefqBOfS8SdBeb0T
y4tddiO1HskqXj5Gl62APdYZ8H6eQ5ZA9vNZamizli5RGXT5mSLNPcPTnAAd5Se2
ivydMk5BpizqE1uaG0i+NfysxrTrulkFlzeOapIywK/Lgvr+nBZEOUQKXZCOaO99
0ddIRcBtftEC6Jw2qQd9JQwLR++S6KoADZnlm3tvEJBELymBDia1io1qXT9dasDn
FE2n9nuV1LfcfB1XXbFVblLsxTFPaMBTHK84g0dWoguSB+nCJyQpdPkz+DvsQads
9V8xN1ICcGcxT5FWWBHe+wusfYloawt3J4JxhZsO44jWtAJDUdcvd9aLjF5OYzf+
yykRfG+Jl4Ri4rUwxGRuDBj86IuaN01TFvFIo4MuAow9A9jatCA5dNFrXFGjOWZe
O2SU4p6/3GeRTb64zX+/BBEhxA4iEnBqkmh4xwpK/lZy6Dg1f88inqTAN58Y4zi4
daeydFVwyL6f+YflneIu+93W2TF6SzwybogVgaiQdX+fSuFi/Si8R8SFREToXA5c
NOzstpn1thLTc0ZiPfOZ5OtTwoQHW1gauMbstsOJL0XwiyjxBY4ryXiwYi8yVDPH
bjZkju6x8CfMhRrMeCP4qmzvoYNPdWs9Y/wG2GI/aYVqBoj1bRTkDEnqaWQEH4GM
WqNngfHCU6UPodC2Rvt65brO8f7MQYqd7b0iOX8aQIfMDcSArlBs9FBQkeH+NXXq
6qUC3z4ViXcQJvFoWoDlJBIchMrDCLSS7sCDMkY59gbcgBibOBkl/ugR/ZlgFZ2S
DOxrXaLYXYRjdPPF2I3HYRfANN7qzuknKFpW8lfmRt4eq4Xl4ff3EPZssFyAgcw+
Qh47yshAjUU4iNbEt8/Wdh7l/rdPh0fHn5+L2KOTDsPBlk9207OOjYvjjtCNO1gN
F8XI6iGiCcMWDeNFPzDiL5Q8hTKR3IdNdYOJsBktNc3Ua65/GJgok/+KHE06OhB9
q82WE49mXvS54ErNu0lEu6qIJyOQOn4JLccz8MC4N47kWYYvHD+Im5t/S+gfEj4f
0hJM0tYT5ODNn8LGdkGWzK4RN3ZlKhaMRFb4Lutye4EeHiKfMMBWNWz0fDTiNvBN
IBmjVsNhwbz1VOT9YC8uKsR8tRZNxSztnnEnrZv+jSk8d8E1Qe0qe1VjlfBvVJuo
669xPgUWYt4V/FvFuaw3U7KVvQUu6LpZHSre1aZig3AAl9qsnuVHP2JIHA8TSVLH
EirtxpiUwXg0/bxlqrXuC+kGNyNcY1/SnzA0uIJZvhLFda85O6fA+8/6g4bq/o43
Js134QLz9SDTU/En0FRAKZWFYiXZUmWzB+wNdmyNEFoGA0Mlb3O6DHwgu1Tgv95z
2w/hH9vUXSc0GrvaG48995P47IQQVxG+2SmwM7qwLTG4SfG9fyxonORTCm7WueB8
ceggr1m0bOsfd/Tmc7tbTIdJCPbZ/5/Q7TSkx0bdsE0Tl56rvpZ3We6CB9qq6jnC
Zr06x0onFUAtKhfjtS5slMNMO+FDt3kXvPsnAT/YVD0/BCGxOb8rpHJ3775StRH9
EG+0sNZxc2jcN6TfehN8JgEKmoDE7f5VhINFBv8fAaHQ2eKjAG4W9fqgs0ywPFkg
BcyEDCQHGeRb39tEhQ1L9JqKmUIJ56/HzUZkKLbzxxW+r/zDN4CwaZ1LJrES7A5F
CVt8X6aWhb0fHA5+yw4yhggopi/p+9pOVEpU+07DWf7J/IVBo8Z3vk72uWNEIiyL
`pragma protect end_protected
`include "xaxi4_slave_emb_func.sv" 
`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="galaxsim"
`pragma protect encrypt_agent_info="https://www.x-epic.com"
`pragma protect key_keyowner="x-epic"
`pragma protect key_keyname="rsa-key1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
cPZNsXIB5S8lusZoX95Xq1Bwyyq350wBiPRWY4NxdAxGbL0aRl+jXM6FcGdXWo9H
0pX0W8vJXwQipsMw9xPU49NUAzuV89tLw3b/ZbMEOdMQKrlOka12CDTDyeya1slI
btlJ87NZr4gZo3E8t2weplUn9kUm7kGGla24gcHQVsfUyCL8U75hFLHNbGCGV5EH
LJl7lnJ8wlvcznL+eDBYJJtdioX4tly9BjCsnL5PruSE5RADWiopaCGn2k3K/J6M
9wjQXNHGmZMIXtRuGmYu1H7d34Ybim+UpRIfz8o3LaqQGB9XhE4BkIuNqmn+3PZX
ceQtEdPab645JSIz5wiI3Q==
`pragma protect key_keyowner="Xilinx"
`pragma protect key_keyname="xilinxt_2019_02"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
Kmjw9dd/3c14r3PELK46p7Z/rm77nhCRv+vkMNcCeiLiBA+LR4gsrqqjPNt2dHsj
zgNUN3skrSion3EBZVmBfAnq4ta8rhCXRuxgUkLbwCo66axInP/zHkOXyvDOukBg
kQxUg00+yDNrY8YOjJAN3qRSg0ObzZ5s6bUx1KUietymk6JOT+TSshpeA/oG1VJu
p5wRjeZqhTf2E3PtS4YD/LQYNf28mTpVfB4mvmZ/QR3Kcu/uD3lSsOvqgxD8P51a
yW0C5STSM+F3fO2ti33ZQYsQnqzQS969kInxDtHIQ+z9qdIaWBQWB199qe7SMU6C
bZs5hUC1CdPh1PGjlvABRQ==
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`pragma protect key_block
qCCDB/hY9V/CNAuz49oh9F1SzV49MZhNwCww36udPNt7+jtyAZzl5dsh3yVzh8zC
hUGjiLVmI2nAwIke3Q8yyf6Si78spr49S2jfMzvQ05uqFfRVbiyYYHva0yRhSHbU
R+97CGYgIWDZlKdZVYUxxj1XVTHRQlwiRGlKz3bWYL8=
`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
mqrINYAz8CNKv5q6awpGBaW9wvi2CQgRP/8Rscx5Xcovm0zD1en5Hi3GSOz76E43
zZacSPix8pFGutJYe92u/cxaSaO2c5t0QVMZYLWv5ekRKc9nq/D2c2Wny+M5xwP1
ncCVuRjbG3SBdqTUWxlW13f4ADXzcJ7z0TmO37SnvXXPCzsUivBWAANSBRMg0xLs
zaTIuJivpYoKngtWaTLbg2xm2RHiX2nWT0b1ZaNIH8nTIJlei5e4+RApHP7C16Ed
bsVo/eWnN3Jd+KIW4cEwt5Yf3ig0G97fQlgnJLZSdqc4zZeBAcBFinx1HxyCxeDb
RMh4j7QYWvizwidroBD5EA==
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP15_1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
yqOQNkwu5vkN5hU6P9M1nX0fnkgfnxjBpiHyZjFD7ZxwCy2mcmtGoB+g4eQnLpcw
3BmsOV1G9soPDYfIk5G1emlTr6Am5qURYvclBbdsR6zdNNq8kALGKzINeZ2sITt2
KhwReRQLWsOgb5dJBy6hMMqH2DVXkN8VsZcvEpaFQQNXKIspfX2jcokc9kVWU3JY
MbUEv9NzjtGVzJVxHJRkK6c9QDlS/9O4zzuAKPvSKeJ3+9BxMBgfs2acalQJEonF
BZs6wddKITt+jrM5YND9OcLwzchXWcjyEtFrE/JZpN/Qen5qLshAX3piW5qyklZ3
QZpiiT0Fe0k9aXB/Rb7Azg==

`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 4976)
`pragma protect data_block
KCPYJh1S9Uy8jB/afSWNsXBzd0EZlunkcl717kI4mHvSN0FznkrOE7j3TWxEltX3
EIir1Bq7kSMyOHkVKpYBzgtU1tGaPyt154Y6KAR0FjnTrJyE11C9KPv5WrGC/JJB
UIil5Qo0fBY2sL/4D9arru9duth/BTWfV8BzuVL5wGovpNGkdnBk4PRNHMBOCanG
6tCtqHY4SR/K2LCeMAc81vHgW/7YPIdTn6OhK0v7/vpAC+9qgsZphHdHD94cz5GA
P0DCdiffT96esYen8IV1hJwOUAN4VlJkR5TaGZvhkkz1qwBpWJ1/csBD7/o93ocY
a89ZOU3AEwBo5An3jWjZDPa6unm5FtqG8dRyxqxU6RoE0YyzE11Tx5Xt13DiZ/ur
RJTbjuYCBaLnfzAONSm27PbKZFhE5UXZkv+zPlNDgp1MwnI3rLKTjEu2dLqOP7R/
kFVcBja77YEyoOkRtv74TFLOcbYCzakC3SSw5B4W4mfZDrGfE6hwCcI+TTbJsQmx
f0q7riglB6FrdZlCBicxzJ+pDjbuPjnOV9RXhoF00lYTFsFM2b2/Qc3BDe2YbjGb
FgA4X3n9grRExANuo7B4T20Ry5Fn8o2jVyG99c+DyNeJ+05Gfsi2zixXfX2cfR1z
6BzGjuPOX2iHEixc0o2yWu9DLuk+X5ia5tYaGmj0gaL27jJESIQgGM/xA75P6Cd5
8dCyZwR8kNqemT/wB9F2LXKXe1sCCHT6IpuPhM95tYjCCoYsJ3kTBCv6cW66hUyf
U+HysyFtCImBUZ7mtaB+oS0faTRyjy4iBGmnzIWRI46uN5DE+I1lNkHFQCy4ujJF
cbr8W9I0V5sezdt1Wu5duChoutbytvOP34jp/iKWEbvG3E7epdewUExutF4Hb9yH
623rs4Ow/ya4eoXsWtoHlEoYXbLpopP80WMcNKPRY2fiRW2XreG24jO+nUPM+WP+
FjHp1Y6tFe23yVLSfsoe6XEs7+U1c5slA7zx4trxLKf7KcbtH+mUvxJtvSOV1G8Z
lRf/PzBgMn5kaEMllEG0Jxy307hX2ulQ8Jp/WKJjThRIyW8gV8I+HvP4YvIMXSdt
LHrYUES1HVQySqCJqeYq9nVfV8qQ44ndb51GzXH1YIScVimXVc7ZO5CmOtyUQ2YW
2Tfj5bq6OFPduQ0c+tjrgAoJbUiyrF5r9NWLm74XcvXQmz0BlBc8jyhcL6Em+JGC
0+W5hQZryn4W3prY0Swia4nhyqLRTFhxY6icJFh4F4Ap7bcNqOp4Mz3+ctlc4DpJ
RGWwnA9HsCoz6XtT1EAim3IbAxRITDeemYIpj/Q6XmokQ9kdPMnNrtU9VB8RU6QY
lRq8dtLvkD0a3OBwOncXIA5LqVF8MBfAhN1GzyGT/2tknt9qVzQKtMrD281RJYC3
bZeAAKopq3typBZDK38WLNCTNeJTMtF7mLlZoBn/V3e9jWoyJRsw1stXA8gIFMGD
n6yzA0SEph5CSiAtts2hsHIejNGYSHFF8Pkuqrw43Q4HIc7449mFFGclEi9zQpoy
YPwiXDFipjiAmRmDDfNs+WHtrJ4Hu7MkDGkt7re/w+kFaNT5gTwf7MHhRigDifd+
3EyHbTf8co0LxbwABHWZH1GrU+WRWAQ/K6WgGtghVda9LTVrBWnoq4OHfeSJEvTS
goDJsF2//WiLVGP2YlXdl585LBrEoz2KKACdkcMJF6UQuwN0Q7xAhdVQfKFZhFHH
4EYweW/RTOebFAV2/3FHL2U2frGzpfN+axmMUX6iueukM7zV6hUPB528dnhoXVIA
iBoa+ZZ40oZAcGHDpQrgit6YJ7q+fuzKMg2tIKAIk4GuhNwadUIys9kcMNB7qvfM
h6qMz9ph5kqv3XL8s9YHckaorfzRiP4xU+IIaEpC9ErMts2qVaRXCPQRKOxCVoMg
rxPrwZh6zmV8aNWhkF2g3UAyqxJ+YR9OrGqQ0zHL8vSxGujF5FR3kBoqM5GGWAt+
zKSY5PZSltyhyMa+gtX1OHWqrN0DZZUAGS+DEmGn1vU2Q7PFQoILaHZ5jxd6ud1f
MIQT/1hDv6MkXcVxcLizXG8NaR6ljmw5+1ZgRNkR0KqqFcaVZdnBdYqb9cnrv7r+
rn6bazHZ0DIs5qkcgl7zMLQQNGxXPngCUl+9qFeMo+cGrm0n77H0XmalbP6mfRfy
RDVd8oPubXGNyTgnLyzASmFLZvQVzPXa4AyAe0l380bzCyS6KyHrA7dL4QXOT7dC
9tvb7+Lc+BVWG0bz98INs1NfJ4bG/yfck8dHZBaD7xNl3UF4W6pTsc3g+ByS8Vfu
oLrNhczGTXL1Umuv1WtzwgcxRsB4ujzk4DtWNoFkRJs8pc1COiHjXqoQAGf6i0N3
J7bpyz4Psoj0JXKL6OUuURV2zm4mYlSrqUirFrgAgIMBYgn357cWyXHs5d+4VEHK
RBGM86Y8wQ2KKJhivtiEavZKZXgNZAg12cQ33rbRIay7bJ7AqMr8tMsJ/981ho1E
EvIOgpV9Ty6IB1+ak8MwvdfHW0rbgwWH9Y1pb5dPuU3tbwFMImYcV0aclswwZYBJ
Wnmgljv0CJy7Kbx5IsGkgU7Mw/I83khBSWqGKbulX/esqN/xStlDq+kvb/ZaC7vD
DZeUAPbEzKdR2B8a2enj03W+r9xBUa6fDsMeCBlB0sdsZ1NwC6OuU61382MH4uIQ
wvshMaoUstqEP+/nVsyb6rCRlssdaCx5kFMaBifbRlhHeDrvdsrmSnlu5F55mzXq
aKbcSENhV7GbhDEtQj+cudgfyYFGZgyCHmJcC2ktAbEiex77ctmOMv7X3PjhOZaA
FqJPxiEXwQcaMkN8uA4R3TSGtlsI29DwfcIY+BN7AKeAEwDkiKRvhC3Xf6Fr4/Oy
8yw8pUp4n0ynyzLmjxYrWoXCYap4/MjAHeRPmGPhS7w9AOkPhqjybanNZZVs6aAw
hjoJ9xggqLDAUOdeYsRQZ5aY5UehpOXV49ydMjqTm9Yk3l5/AaTBWVDDTrngXHvs
HmkqREaoYwFgwE5y9/1JiBKhcHLIdOP76SxkZIYMB9PaxQ1o39y5qZdESJC5k8tk
ng2eYi+jJVpaZGfxXx/+X4aTApo00WwW16csP4UahSoTdIUGK56AgChGfuniTjUO
67Qz+QXWaXhIF65DA8IXlOVTUnoO9dK8yuLrjmntiECW0Klv4mHVyTxTrZ+/FMog
1OGHkmPAjQl6JkEoLyOpPIeCwemXYcTfbvkAUi/1tmQyx3tfoiIlTMNwu8fK4XlT
mx9HwkkI3Z574S9Ddp3/YgHs4y5geVDt43P6zGRQFMh6QNq5IcrOgiJmEcb5dwp+
9bOfR/QGFZEuN4XzZ9b4fEERedNLlP+ftVHZ/HqYMg60ALfpx/SvHRKYJi0q7zss
UWDzfvsJZ6hXvz7pR9Hi3QeW8sJuuz1UneqgwiyDfq63lYSk8V364uZNZoHx4Ocy
W38EL43nx+0v3w+wRMJILexUTbh730UVIVZ6Hbh+Va74PHQf6hUooFYqz5VIChT9
htk/8rXp8wIFAf2/+6DkEvofCDIezS1Ni50SG3qtqLTQorf+orax1f7bDuJI+mOi
XaAeJ0QC5HEF6lpx8uR0OO1b+Z4WAxhBIahTazxCvHTVseSmquoJSxtS6Z3VGDAC
KgfdT9oaGnpHhGHMRRVhX7jCc6Z4KMrKbMGDNkoUqDRqSCFA8JWoeWMeUSQJICz9
olUUUPrxs2+wzeVa391Kfkd4CBMkn8SiW9/zngSX63JHjAQ3VV6MTDenox4roIy1
xCvVsF3f1geClVGyuPHvoZI7f5IotW9TCzbRHwAT56Re7muECv37+WMZwmDlSRcv
qlNd4e9H8/piRxwGU3aQ06eXbd43CJ6Ca4Ss+x0NLPJhEMyG/k+WsbPHygMwCxOH
p6ViBSAsZ0MMeoqZqpFykyyOT4Pe6IgtfmKRPTwts5+W4OGSvuOx3k8q0hNFExmJ
kkekLp4em7ncvmImoic0z4zCbjjzGUSpZ35xw4b/FnpkyIbhthRhIECCAlTlqu5h
iuxkLptcLnMRDD/o1kj71WZaysW6YK2U2EEMlgHSnXp0XQf1m93QMQT38d8THGC/
dp870yk4MbzSctYk+aTjH6Rv80wTxxvAfMPSgZZqM8uL1E3eQ5fuwSovrEFFYh61
TaMf7jV7YhRDc4Jzrwsl5Jd0ckTPmmSPalqdH33hCzXKDvNzxy9RcbrqLCNlTQYO
1/TmTasz9NiV3WY5o/qptA54/uHkzhcF7J6TdJqjZl7vK9Gl6GWtsf1S2hRXI84M
AXS2Cc/OGWQlpPqF5K67zeZjzmRLIOKk/pHBCRULNqvWFmZVrpCLFQ+lvVIALevW
7f5Czd1l6GaTPsly4sDrF7QpUDRZMCHB9S+KJKqHDx618NvkhSpEMuEtM/piUjam
oDcEZkeiPPLwfNWAouifk0uHY0oNAe8iC9fbwpXrBwaudWKcsisGJ5vTUG+3g7Mn
1lELC48HyzBoxLIpF3XBRUp+0NCDT6ywcLbFKjSEuLhVb3QPvYiRB688tsYdE601
YoaijDCZy05R3Y7VlQdRvO6gThiv5BXjpwpLzTimLT0epLz/oGEcOYuZmunc26yH
HxH1bhQzY6NX9RWYY0psbqb3yKwjCCTfpEs0IZ7lrwhQcKOWW96i8wzMc09HW61e
2o6e37ajrDuqQnRA+UIkItsP4WxvVehU0kDVBbNVQGWZl1jDp4RtH+D0IVaIYZX9
mbW7Qs8DUfaYtikxGdKy6psjgbZfJvnqxOHhKymETllc4JCToa7WHevt4NYNYzE4
xqqQedn6GBpoh5hn3OTgScog3DEGtVGtRca0k+Q1TdJZ1IZchEBL3mRhxhrIf11D
zqyWXaK5W3Og8PPANyhLg/+joCYEawSy/qF9Uxav48nWialAmQyv5c8dNa3KTI+3
QRNHlrWSBG3+NCA866FiIalzEnr1pc9yL4QiGAY+4rofLDPqCvVZu1qoT7Pxgxu1
ac2mN0ZwkJ5tDTLgjyKDYVJl4c5lt3rPyOMk9oY/5kW/g0kzOXhWdgP7c0D3M0sF
+UBlLsx8w8nq8qV+UIn4KXvLB4BRUeTNfetmKVbgsHwcaFJvjAcaN/Ooqy4ymLIJ
LytwizkiVl9zuIpw87njErdTNqc4Qv/aOGeTY8v7FuJ+jvh8Jeg+qeyoiHnp5pcv
nEl8K7DdRrr+4nPJG+tVFcLlddtrKXd2kAvQYTMDeMGXPY0Hm2u/CoTECJEagVwr
3CPTs4SS/DrpicGRl/ftGYpom0RzG5mHWnc6kN5zujzNukg3ijPKDM2tOCLfMREN
//kVc+MULiKYme90WFX4SuX9loU/2Ny5RZOwNCxa9XyMeoD0Slv94gqlCpCzHSSz
TieACYx5AG8eEM9uHQX6w2EG6D343lEXgWdJQ7e639RPYQdWGST/Uw7Zl+xL2ixU
W1rz0jxMiLuhUN4hl5bswwkA2M7noJ7mcWKy8lx9yk7GnUddV9bp6Oc2w/qL13dU
lpqzluTn1qw1YtC3Tw49TJeLOj1A3hHOGvdfw2SKQWeBodMfeWN0aVgwoyOOHbUT
KF6hKaeGi/KCU/WVHxlQD80pXi7VPKVmlonEfLG0T7vFfLOTfti9XbuOGG8Twvbh
6QOEl0FgHK49kKp2G3vKS6GC4Nr09LtOeecKRKn1tRIU6gC3BztT+2JduAtk3uwN
9w4QsyNkCg9EArN4P8waYtVsiRHmRIefcCeoVW9e0RwTyf7sPkGHSBAos4EdlMfT
vm04qCMdzU2TypcFNaQu/DjGXi1fIiPkG1mhlgJ6lyjqXB4X3Azs96D2cKKoRr/f
mrFT/82iMBZEzuuFg2Qbwz6Zq1DmwGIP5jEtEAESKWzaqmn/IOoAoYEEbAVVK5J5
CvJU4EiKU4Tcx29kG5+drWb7zmqKMZo/uapPad0SdsSvdbp32vfRlK6PnpqMizzp
yBzraV6BLyeE5ssuVBA5ZS/N/GuACayrsevZMeaJraXLC67jAQBezerVAYORHmb6
iU79SEWxr6IUA1S5F5BEAy0zwJ+UMPi5SH8OhL9ZoCxMyD9QNhJgNSOp56s0uZ1u
lt4mFNFN44lLZ6a+3tB2TyLaU930RXKtcngjc2nJbjxFHW2qbdvWGTgaWwoVoMvP
HJitm1WGTdcFeKm3GCC5e08jnM7aV60+wkvTJ6dnTLeepELLiKw0EpXymZaRDCm1
JJt5E3W11cu0pAffE7CPo95hpMeo5pG9/SVo8E7PcNsnqGMgJUH1wYMvnu7qNvyF
qV7PI/iPYm0vlwRAAq8pcAgQCxYiBvc+HbAVZeMxeFDVsCZA5/aoNmjL8I1+tYV3
4NXT4k+7rgXXc6m2k2yF+EMpKgFdMWiv93xz3JJ/VtJGR48kFcnnT9DP2Gr/oPu+
VvFeAlaNf+RueZNNq8cWJHhIZXCVA+Ju7s2fxKAB1nen9Ry9QEZbFBOpkbNMzPXc
IQsw2x6YtbJvZq14xb0u49KTbkyulUlu7WSkVa9NMlNoeD8CqIdBKVm5nH7mi513
vBRPYhnUwsVqIzcUTbmW6Yv5Cpba4YkJ5xx0Z/OMzi3kynRSVqvc02p0RmAjQHqH
k0okiDjgQvqfo4p9g67qtxlwA8UONnPGElMghVVXwOI=
`pragma protect end_protected
