`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="galaxsim"
`pragma protect encrypt_agent_info="https://www.x-epic.com"
`pragma protect key_keyowner="x-epic"
`pragma protect key_keyname="rsa-key1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
jqeH6nkRk9EAxSTl69764/ZQ3dMFfE9RUR8At/iKbt3NqXtf5Dle/EotUGE0Vyxz
cyiMydNgVfCzBAJuB3Fr7jagR4p2SgR/WUuEcUFdkf5nczP8dqDnUJDk/xcWnMOV
PosioXNuMLf2kD67AwPmdussP3tCV5DyY4DbykodKWTh2IqH4Tnn5RunaIGu+2UJ
4HhjAOHYO4j6FMmxXzLjlyEaM0jenJNFuUR1peJUTnPrCnVcnf4jL/ZmNzRb8p0j
93zcB37t+EvwRfcvZfqz7G4ys6dGzD7tNqHSgfnJrJQwcwL1j3KSulUgOqm5XJ+S
vmOpHinqDwGES0Ec6RmsxQ==
`pragma protect key_keyowner="Xilinx"
`pragma protect key_keyname="xilinxt_2019_02"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
RBpx98Of65sgrGJlYgBTgs9sPnvHk5lVIUtNRFqI8kcsS6sSatedPY7wrRWqCTuq
YvoSxspFSZyJJYkgvcFA8FB9nQ1YoCKnIOs4wMEg68Wuj1Z8q7k4zXbv1+dfd/NK
C4LErDe6Y2fgskMbuJyR4kkU0sB0DSB3jwHpLNMkve4NlqO4VrJhyHtUfwFZHhyP
QtBNGuHyMjDaSZTAXSD5+hxreL3NV36Z4VDpShxcsDfAXpdra853S25byzfR8Fp+
5iF/1wU1WK1KW0F2IGBjQ/BbTb5rxvO2qVSZ0sLPK3goRGedt/7TZoj+06EgaJru
hRe4/QIn78Td9g10gdlhRw==
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`pragma protect key_block
QJmXkVENAImybOz/uOtOeehNo3OAwuEovYWv4xxabNWQMs5NMriD6v+VMlaK+0Ft
VeQghsauIsW50RkM1WewfFAYGOtltaTwCxUrNbiCpT7lyd99Gu36fZ0UUimab4pn
n3CK//I8piBjTw5RMBK6r3CjpiSpoZXitwO+/W5yn5k=
`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
UEeY5gGhIrWq4RkMkimID2YAabBBhytWqOGmltCw62l+Ti+wDVbHm65a+p5bio6T
dzvMFiC76RXWDL1OMjbJ+SA/wo2G+HJG073Vlzq/oLAxCOqSiCxinNyY7zjKrmlI
pynTPDYbH+hEUM+SjNPyy9599oOvqXEXE2fqMiRLOwBVmk/GYkMtpazEJdoJDplf
6vBfB/MID2ioVs+LGN8IS43SRivjmgEwSKroOlCOMkvzKziAYL91zQG5XqMrUhh3
QS7+zZ+VHF0G4pgyZuB7baLQCZ3voA7pSi//218lT1Jjvc4MoOlUnpWUrPiiULTe
DCA65FXiqtm+8UT0i3wZDA==
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP15_1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
bSJfd9JffxjyklSlmGEEGlWQiUESzHg+0foElLZpSjlmWFJzIWxL7b/6r6kcVAEH
qxr7dSDV71Lmea7SOJdAax8fdDBAmYBBI3DkDPj3ObLzebLXmPre/BLEyPm+Z90l
23ofvmXsS/BxLxVJHlsISKBQ0LrMOkoclyqmRJuoCfQVzNFLw7h+KfIo9ASYkRL2
NB1tFRaMMtMEBkzsPt428ry0Ct68CHsugTE6R9jRRE9O4U7+qsjAdHeqo0J/YUJn
U3yEi+1lmc/lOLAWJXxkNPHT6oW/y+pOKG8d7+muRY/ISL1xVsToiD1Y84kdLx0N
rp534OW1BRwJbUduvxRLwg==

`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 816)
`pragma protect data_block
XzAC4OsUhRVi123o2eibwRsYhViM40wcsX1NHzoLq92Mv42dflZW0Br0MRYD3lkF
q3ioAg7T9UrpGTbZP3mBLSDVKcRMTKv/SpvhScALIRkw687mpN12UxkZKaU7uyjx
07Mn78a1bS7lWgU/z89zINl0S7nWlAWiTDYpxi+n2Z5oWABnVS7K9lI49oeuhpEk
DRv0ZRRqKeYFQU9y9NN8EJhTCxBcX8p8Kd0NH1cqrtqTE4bJxUb/3J/Lj3LkLkYz
7DwRUyrvi9kJ89pk2R4wL8iJ9Vp9NWoxSokDxqdPpMTLEcHO8Gj1Z7uPjaJR20t7
5FhS3coRtHg1NKgVO8in0xaaPuENJYlCrJ5gkOtW1jtumfWkbUuw3OTwkxHsz/Vl
t3AUxQz+e7wZJorm+aSt+PhLxROmJFJ5sIiJvYp4Ci/2rIrqEOIFk/0dng4BG/Hi
AHCiRoH/e2NiFsTVzr/56m/tU2nuHBlIArF9N4L/AHfo53XEnSfXrgICjzbRM7A9
fDMYyAsXWYp7Y0ucRhzAS73tKjS9x4dNgxzGXcGmfhtS7MgyTIMHCYbKtclK3nGn
HxAV5EAdZlyW7iRp1Emn4S+hXBYvrnf0tBGbI1I0CtbeJumEHcr9Qmefpcm98QuV
apDfgUtal8o292XqSfYg9yO2yImaTtLww4iRvKdVVC5e/7x9aoAPeQ1jXxc3agZs
Vm5SfJxIFFrW9upfO/MwI734taOVcZCIDw4m852ap2qW1yvnXCDanozuCWRohJcy
UeBBAyhPd0AXfVPqEdeBAzypcS7F64Ag8AKLSeD5QjCts17VHF3m77aVQfHgiicX
bt7cxkS1aw8waYj/belHa+tIZ5JOvIqGytBs++Ya80N68QQLz41tphl1HsXD/16w
tKkMbj6B484KmG/44VD/+xIal5AQBzsBOQAjXDJD3+FsUy3DdQow0FgTwonTmaBb
kn5cpLlMsa6JfjrJjx4PIxpXmHGwYn2PJyhv60r/hgTOHny+B9XeT5e7PdKDBMjP
SAwG097yAEc+wKcfZaHWHeK+Pb1T5VqjdXkRd86SQ0tgJmKQkm1KTsce1lNvCMWd
`pragma protect end_protected
