`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="galaxsim"
`pragma protect encrypt_agent_info="https://www.x-epic.com"
`pragma protect key_keyowner="x-epic"
`pragma protect key_keyname="rsa-key1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
1IJoxM2IeYJQtTe/nJfbn41RCpo9OIxljK+YCofT8vm05ojiyu9XNV146pCdA0Y6
fMCpD4MJEJGDD+QXKQomj8gKEq0QBRS7hxF15TDB+JLb4EjAa4OIcqR/Nt2iWyHj
glBeyeCriur5qrpyWdw1gjtvThVEMQ+3ADVvJpgFL/YWV6GY3tNhQa1QZf6SFVAn
zzsdf/4N6IEAjhEjHyYrTAflOAkS2Bv8m1UekH4MIx+RCA6VfX0fug7DjCiJ1vuk
D8eBPvo3TlfX7M2gIJWqBiogWgeemzwQV0IqaD/El7Hp1OAXYKnB/Y7HbFUX0hV2
ELEyocQtzUQEJDJxVhe3mA==
`pragma protect key_keyowner="Xilinx"
`pragma protect key_keyname="xilinxt_2019_02"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
h0li3JfzshPGMroS50uNjD6wuTvXVzt91Ma2g/vgzB/0/a2fEpm071vgxnOpUzwr
KN0X/SDP9Oa1BZYB6oOW0+5XcYBrRG34xZ2QBwxx+x+mFJ/Z20Vjk+0hfYQ8KBfb
JnISeUB2Bn0vINurBiyCLQ9SQXDMypsij4wAaQs+FIKpLweLYB/6GCWTmSaw63i0
A48QSoc3m7Yyv/uSfsqcIC3hSlip5br3QZJGiTo4N+aV6LF5lM8yJEsP1UubA98y
oHqeO/7PPKU6YqK1mivPExWxOlad4S9NCKsrJ79FIN3WFRWRoa1KJqHeZypjh3Rf
19v+ptW9PZBkFkRm92DhMg==
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`pragma protect key_block
rTldS+uvLYZvRtlaoKP3daiy9htkIRlluaGOGTUTSMvgj1TU/+X0gqGUZcdHZDtc
gcoBzMyfDCRzFlHy1noPEfYJ0M0rK74KIPBlujedQF4x5ppDm24f1UrspWJ2BQcZ
aYBZ5aCFQzZckaP0a9joALjJXRPfb964dU7lULanHfk=
`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
XZkzAh/nqfcaG1FmCSe0MShJrQN8YGiRwC+hokqeynzakRNkPLWKo4VD66B9uZIC
T+CxfaLDYQLcpirYC7pHYBGHCL4k+UAj4T6D1BrTDL2xF7vWry3dsY7cYjlfSI5+
xFtR4Nu3hjh9WW5r9v1DWPY/zXv3sL9I8HX89cnIixXd0YamjOlTutv304i+XFRX
3V0DhX5jCpSYmTUiW4McTm8EScOHCABrDNdj2t1OjsQ9w1a9uuolrFTMXGx5JtwT
8R+RZh0TRJU3Ea4pGqAyjGjIlYl3QHkNJVKU67a9f0wc7sbb+d11ZJFGmXUaCXKH
7aBrEY17GJi+DGla5XYrog==
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP15_1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
JaEQ+nFmwYj3gRODFHX0Si8NMxYCSTszi8ZXmm0uwg84ts8lrXH/AzOuQK+M6vHD
j6EV8jU7BDUNTtH6PBD1DmNK9Ohd4JFz1ZqgxxY1yw+O0YZyn916eM1+BoOy48bL
Ezqivdrspc2O4ySZYIofhR1pUF3nS+oTAIOsXO5pAsF1VxTmOI4irdR8U0RuC0rU
2OLFx95GbXfkEbvwbzpA90rktspIKC00JH4ElexFrP1sp1Rl6C5QQaZThTJbsYe3
jcg5EzNhbxzrW50jUmWwl01Ixk9kGA/7RZ4lzK3adT67FX8mcTBaGcFfV/+xZa3h
Radrwaa0ezuxH4SxVY+yWw==

`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 416)
`pragma protect data_block
Y+A3Fsouab5IA+7i5Zc1azeDBZR5Z/A/XiItS9zQiGLD1sdKt6TILiwjaMzLG6OR
4/nsCTDd6hBBkG/woeGkfG7gFkMLXZWss34GAXOPoAaAtpF890jBNONPFFOdU3Fv
hKUyHrRNkQnL7teQwdw9u2Qf3tgITTxE0apBhHNMFLdFIf2+P0n4Gz+ahriB+DRC
1RoUWDjR+LYL4UFOW8g3ziZMnL/wJ6yaP2T1ko2lytBZHsOAz8Kfixbq/PnebjVj
jWfhGcdv//kpBw+7+p/5hohyeHB1HSRmuWqpE8T444ic4jMXU4oQJu+ZWp3hD5d8
Etcy3or183Hs0uQzS7LrzNvX/4iy0/MlGHalDOc6F8ayrCHapaNhNCqnYPfZYIS9
MC38q6gAxrTWvaDh930h6tz1oA9HTJ3bp4LzYhE1NTL3pJNVpLJDRW97IRYJs5LM
ZtbV3oO/QWvDboCj5tT2ZyXE+3vjlXR3XfGzsyIpWPDKjFRcHaumckjO4eGzLbD7
pM4LGjFb4/bkFTXJsqs8PyFgCMq5t4uWu57WM2qFXr4=
`pragma protect end_protected
