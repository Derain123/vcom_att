`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="galaxsim"
`pragma protect encrypt_agent_info="https://www.x-epic.com"
`pragma protect key_keyowner="x-epic"
`pragma protect key_keyname="rsa-key1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
MF5IFIGeWF/+BAiTtGnJVFJsfMzpKnrLMdGJfZU8a1plWxYky0ykPiSbAaQInX3p
xAQIoZEgeoOzNhlh6VSzWqL9etvfwGPk55dKyfwDEt4CF6mGUR2oPwmsRVmARmMF
t05ZSxSka87+YA/kYJKiB/WOOEzTaF/eAXfnhwnPef14Qv1XVHeGBlpJsED5IyFV
AlNbbAZUZiji9f0Srmd8eDu+yiFyHztnqWmaTc9r7oq4gxWg7KOQkwuT5MIYKZH/
meRvPf4NOq0ZI7nmXf9r6uV58Q7wubnjTFfiiDoKMbQLJ8wZ7T5sbRzAgFgQ+zWA
PVFRUK1OxULtij+Ws0JjrA==
`pragma protect key_keyowner="Xilinx"
`pragma protect key_keyname="xilinxt_2019_02"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
FnMfUsSN7mET1BQQHqmVD1I98HN8t5O9Ei3RqJocbzHKRS/aNhbaIAi35ZUv/Q5d
0844Lc0m5ZlkQa6jHMpy9lDCkdOY+O4D6bQqhm70wsTGj/fJ3sJQt1VMJE9akx2j
DX0OLO+MbGtgspbhMZu6WO/QFeWph3LYPsvS45+j19M+bbiieoh/Dzee8jDcULsk
Fn2yflec08aS16NzWHGXVoT/Ah3Zi2H8mF3c1NKzig8fjnP/wJy6aYgNAfBsD1OI
sIb6S5eaa/dAW7r080yDHHmXVeYpWqA7qTTDKoJHxuc0vv8k3ceJJrH+3ZIt64fw
8AIrJBWXJ1w/ekV37PZ4Ng==
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`pragma protect key_block
Ut6unzHJahSyeXuZCGIJAgc6IpwTQWQOK8adNJukFjycNHmhYJC1dDd61x1MlbAO
rq465LCjuLZdkftEZZF8vO/hWPlQUs83IvbQpAKDZ5KkwnB4XKQK/3EIHTxaCvFa
d4Os5za/lw3zq/1OxcMlV8gkFFfNfrmFdYlUBUagNgI=
`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
p5FS7/HepGCSyfpXRhqJQ1X9lScrJ9DNtcFjhJgf0gOrseSSZtC8x/AW96Bc9C2W
BYO1sOSFtm+5Kl0o+lnhQb5XsOMupLM4bMeUGIGrDJ8Q0mt3ogSLS72JTujNxAfr
QB13bpilonP3mvqoJ7DafosKdHzGb4okGYpKyMb79oTjfc9HbpYuiB+laOdMqM3w
m1iuHOxNlasChpk0TRu03UMt9T+e8DTFus2FMHS08bEZ6H83ASAQWf3wczy09ME9
nvOlh85ZgsrYCCnxCKOg1ldQ6hlX7R2j4tDhJTAcVVtfW5nWsWfRJqMYZs0pla7i
xaJ6FEKjwVA/RLvIhmYFxA==
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP15_1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 256)
`pragma protect key_block
cuwibEWAWiJwWqk3qdfxFpMbXcKxgrINZX4DAbDw1Ff/jDYbRez44bgF7ouPWK/W
hP5VQBCUWLyKj50abqMq3sB7eOIz/8UgccVFDnwa+/LKUhR4aFBWDf/NDXNI0Xpy
HDgqlwDl6thkskKN7rIDIyRbch8ffwXhjW2XCGA2ZbOW2MT7/i1YX2Pz5WDg6jIU
PUCfxDQ530t/mxmKPnrhrCXPS77QY6oEdkUQ91zLzbex4/6EDUik5Mjp/JB4UjjZ
wkdpvkyinDVZ72sqVozrRnAHruZCAfbf4sxVgizBXQXBnpmWYlrWjF4u5jnCdRVi
VoVw1k27q2cTo6xMy6IcSA==

`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 2544)
`pragma protect data_block
XrszLZDNbhsicgTXbiPRx/TCVNPJcZJwPLq5N75FrIxANHDeii9y1g25JgUxywzM
IA42ld19QuanOCEjualnsJK9+/HCUPzi0ye0r6ZW3El1MkvTyS2ZaF4QBbXet2Zp
UPyeXTQcSJVI2nDvSBV5ysnqBt7QEIFXlqamAha4Gwtvv4mpQARj3cT7o77g9zgT
V/lHpUm/wGXO5u3K+Ssn5uaWJLu/FtPnJzVj3Nj3/+U/f4mAdV70ji0a6Eb4l6UH
lqN4yX2a+6XhJ50VtH9G0SJhsPVQYWKQU1LvdGtDGD0M17B9RCbWIZhbvO2rfhIV
5n8LuUCDX+lYkjTuBYrd4yt2Kp8TWL3yoIQ/1r0xvQ36DDnGK9GOv4erXWvYYzaP
+NNBFmLtmp8+Tz8Km4IU5jJhBPzHaaRu+5ZuO57EezE3XUe0stt5FrNDBO4qZNeH
7qShHf8haO+3KfFUoKYjH4AmfMalJU3G+rSBP8dcWG7CkQKD54i9rCxxagFF58rB
FVQM3NPmMtFK4ni+RWctTt1ApUg3o5cBa1c3HHbpW+0GgA9Xt2kKXpPsX6k4xTmg
RL2J25CZeM/htn5pSSQnMfM7ZRMdv9fMZeyEJ/WgVzDD56R5rDzTQqQoWgezKBdA
fBnlYSo/MakjS9LQgml6Vyr8qMul5EjbCb2lgg8iRj5u/i7H+5QxrJhm6i2EgL9r
Bf+116Tm5y7nwYX6phPQ5KkjqR1qeh2dOMhBdwOq+3LnlN7evdlaM6Xrw/Ji1ThX
QNL4jMEmjyhE1AAIitllQ2Ybrti7lXsaH59jcOIVNFRAjQjCaTJRyBUjiHuSkNk8
rd4mFrlYqX81hXZyjw65VKrixdZTYqoZ7rKp5/raCbFiK6SkFfvfzQGQpg+wNgfY
Nu0ekdegnQF+xS8KTRaZ5mQqm+J3VzjNaL81WxMzy7CeE5zVmZQWld/leNpPcz7l
iwJNrp8y5aEqIx5SxDMJk0cNKtlxGLhTdsgMX2kMU5QR3au57FKwF3aEhUobLOCX
EJGakL6FCtMYrhKtM14dytza5S7Qnk2w9KlDxondj7/dZ7C7rIVEzFE4YbI+0WcV
+BUQ/Lerlhu/59CZghwYUjrFHALahpy0286j6Slw3jIYXTndqrQa5h1HiRTwKkLp
FwLtBS9Iv6I5A07rGrN+e9mjMNlTqP+yzuMkG2t8NBZkleP2hsp77JzFQ2wdW9cq
N3SF7r4BN57hJ7NLIPpcfenUSbcr9P6gNdUkJ/OasrPnXf7ss1BL3qpYnhLsnxKn
kpNQgL8m/zsT7NuHypeh/8amegj/GJw8URUa1gzHaU3qmhhPJb13erCPxngcytJA
S4vYzzEZUG+N/CSVF6T8+ozQYno4gNPtisUxMj8R/1Xmud+wI3NDUWLM9Zg1qloV
mKFxV7fwQPrAb2CNxEu90n60DB66iXs6gY2xOUe7wBX3VQmy6Og/rHgjcYz5XrdH
CEtjG9p48O4YfhG00pLSriRZC6FwTjWgO3ggjcGvpi9ddtG74f+l/a70M0Yf4/E1
Acz5CTIYzA0U1cHA71GQhtuqmhE74CNw97T5C0BWmGacVTcImTWp5bAwnz5ZkuGW
gD92P9EBEZpn4aWEgoZ/y8hOshicwLufGx329K9wbWEq5s0Qvw+m8r08ZZ4MWHJh
6lrTlquyJKaimdX5juqOPUVLkiLuctI3Zb9j3xFxCfi1KsicueKsr5How48mQ0e7
m7XMCo/8t1zG834wctAmvefYBBpthb3W4sDcQ1YUmru1xCZwIGssOGUK1BppHc+x
OL2QjC8tPT2ix0fC4XO7dnEPtyGg3NPB3xY5t9TeL9WTfUox6BzfLR5Pvx8GVM7P
mAL+bUNdSdTrXZ2BUDXpW3ueZlaxjevEg4cF/Yhyzt3e/8OwSt7sGT7RwA1OXcYk
gupUPWcP9idQnbArrIR+Bx8/lU/THRsRDTDPBXhKZ/NyrMYgUMmltaYF+HwAUzxO
1ULXmLT2U8agFDzXyyxSBtTKjHlapGxcps0YluYHuulZGAh2Oxk0pxeELe0L34w4
Xwe5O2jwMufcq1ZVFue9H4FS4sCR14HZqGf/+Y76EGep+PUkKPdeaiVReAZ30fqE
ibJrHhhELdFlcJhyDeb++Qpa6Z/FpRjIyrz8ftbZ0vjA6ufD3ugA731W4Z8Mcjer
WiaKMGmpHgtQxv8JD9td5t/m8grKtuGxq2agOd3izBNhliV4E4RCT+idOoOBVOic
ntNoS/po2XSxZRyWDqDxGjwaOULcYVJfSGgSb5X8ZVXFL+8/A4zZVRDcOTV8uhIa
sKPV/CFTwFL4Fpexh1mQm7qNHSv3v0FjsHjcB+U0glPoAJoAAJEavaCdqFFf42HG
aOIEXyXCSrxDpKHaP1KsCn+516evMzbNHsoAyFshgdYIeZWsC77konRWK0qqjmfK
rRDYgjY3eXyaEXvB84+4DUGdHkr/boK/xIoRpbLJLDg800EAcV17IO93W+1fntj9
WM1MWuiM5gx6kDkVjAtLt6pIiYZm91iurvD8Pn6LPQAXXIIBg7scU9yUpVnWLef3
IqLwr3AudpSgFZaZrdryI7gLd+sanVcMvUrKZ/ESrjjYZwJ4cIeepZauxVtoKYSb
4MAm7JzZ6iCT2vWPD0U/8bBxmDvpm0pb0nVJFzE3iQpuVxvSWUqz/tEQA3MydjEs
NFSmTUVOWP40gYA3YeHC+LUCvuKmrWvDAH/kPL0Xn8gmtFB/4iV6PJub/DYFLrAV
PzSIcSPuKV77x7EjzOg8fWvCw5Qtct019xBoqSAF34Gj1fvASWB7GeDsiwCAkhmI
ly8eslzXH3D7m4FtmM1dq52Mv+a/bROCYrL8javy3dtQvV6OBNDOZmTDeqL1+5Wp
g8i7Qr7UUtPTT+o/b71+YrVMbsreDeqAxkWqqM8VasCvDJEGTmTNoZZFGNAIqf82
5OKvAeYMP0KlBIfVbcCGfKvSuuAJEajW9WxDit1O+3pKba3YU1EB23c/bP5d15ez
kttmn+ubeRTEvJcJQqFII2andolS5a4MNyqyE9igwDTaguM1zTtiuO5lJL2EWVWU
q264+SmFb/4hbK17LuxFgXRdNxKhvSP8HBYhAGzqubeqrpdXwzmCi+msaqjEwGgU
WEvfGoZPp9KRQZmtolYPeaIJha1wFLiPmJ/oAANPK6kerdSrtBGW4WtJ2x293v9+
JX6DiuyFjqobnGDv4J14HvLX/gE5iHu3Y++lgAWvQFnc7jauEqk2NzpRhwhjkFrU
+d/uopcxZtFNcRoYCe7MQzAM3XAOFnu26iTiSoVOQzOX8hKiOE3uFjVf/VNc53CF
MMtHd0Vbq3h2WKhl9LXpO+P2qFa+4oVAVa7nvozlwxTkb2X37jLZK3QcFwc89uHu
`pragma protect end_protected
